//Generate the verilog at 2025-08-31T15:02:47 by iSTA.
module ysyx_25030077_top (
clk,
reset,
ALU_carry,
ALU_overflow,
imm,
rd,
ALU_ctrl,
rs1_out,
rs2_out
);

input clk ;
input reset ;
output ALU_carry ;
output ALU_overflow ;
output [31:0] imm ;
output [4:0] rd ;
output [3:0] ALU_ctrl ;
output [31:0] rs1_out ;
output [31:0] rs2_out ;

wire clk ;
wire reset ;
wire ALU_carry ;
wire ALU_overflow ;
wire \imm[0] ;
wire \imm[1] ;
wire \imm[2] ;
wire \imm[3] ;
wire \imm[4] ;
wire \imm[5] ;
wire \imm[6] ;
wire \imm[7] ;
wire \imm[8] ;
wire \imm[9] ;
wire \imm[10] ;
wire \imm[11] ;
wire \imm[12] ;
wire \imm[13] ;
wire \imm[14] ;
wire \imm[15] ;
wire \imm[16] ;
wire \imm[17] ;
wire \imm[18] ;
wire \imm[19] ;
wire \imm[20] ;
wire \imm[21] ;
wire \imm[22] ;
wire \imm[23] ;
wire \imm[24] ;
wire \imm[25] ;
wire \imm[26] ;
wire \imm[27] ;
wire \imm[28] ;
wire \imm[29] ;
wire \imm[30] ;
wire \imm[31] ;
wire \rd[0] ;
wire \rd[1] ;
wire \rd[2] ;
wire \rd[3] ;
wire \rd[4] ;
wire \ALU_ctrl[0] ;
wire \ALU_ctrl[1] ;
wire \ALU_ctrl[2] ;
wire \ALU_ctrl[3] ;
wire \rs1_out[0] ;
wire \rs1_out[1] ;
wire \rs1_out[2] ;
wire \rs1_out[3] ;
wire \rs1_out[4] ;
wire \rs1_out[5] ;
wire \rs1_out[6] ;
wire \rs1_out[7] ;
wire \rs1_out[8] ;
wire \rs1_out[9] ;
wire \rs1_out[10] ;
wire \rs1_out[11] ;
wire \rs1_out[12] ;
wire \rs1_out[13] ;
wire \rs1_out[14] ;
wire \rs1_out[15] ;
wire \rs1_out[16] ;
wire \rs1_out[17] ;
wire \rs1_out[18] ;
wire \rs1_out[19] ;
wire \rs1_out[20] ;
wire \rs1_out[21] ;
wire \rs1_out[22] ;
wire \rs1_out[23] ;
wire \rs1_out[24] ;
wire \rs1_out[25] ;
wire \rs1_out[26] ;
wire \rs1_out[27] ;
wire \rs1_out[28] ;
wire \rs1_out[29] ;
wire \rs1_out[30] ;
wire \rs1_out[31] ;
wire \rs2_out[0] ;
wire \rs2_out[1] ;
wire \rs2_out[2] ;
wire \rs2_out[3] ;
wire \rs2_out[4] ;
wire \rs2_out[5] ;
wire \rs2_out[6] ;
wire \rs2_out[7] ;
wire \rs2_out[8] ;
wire \rs2_out[9] ;
wire \rs2_out[10] ;
wire \rs2_out[11] ;
wire \rs2_out[12] ;
wire \rs2_out[13] ;
wire \rs2_out[14] ;
wire \rs2_out[15] ;
wire \rs2_out[16] ;
wire \rs2_out[17] ;
wire \rs2_out[18] ;
wire \rs2_out[19] ;
wire \rs2_out[20] ;
wire \rs2_out[21] ;
wire \rs2_out[22] ;
wire \rs2_out[23] ;
wire \rs2_out[24] ;
wire \rs2_out[25] ;
wire \rs2_out[26] ;
wire \rs2_out[27] ;
wire \rs2_out[28] ;
wire \rs2_out[29] ;
wire \rs2_out[30] ;
wire \rs2_out[31] ;

assign ALU_carry = ALU_overflow ;
assign ALU_carry = \imm[0] ;
assign ALU_carry = \imm[1] ;
assign ALU_carry = \imm[2] ;
assign ALU_carry = \imm[3] ;
assign ALU_carry = \imm[4] ;
assign ALU_carry = \imm[5] ;
assign ALU_carry = \imm[6] ;
assign ALU_carry = \imm[7] ;
assign ALU_carry = \imm[8] ;
assign ALU_carry = \imm[9] ;
assign ALU_carry = \imm[10] ;
assign ALU_carry = \imm[11] ;
assign ALU_carry = \imm[12] ;
assign ALU_carry = \imm[13] ;
assign ALU_carry = \imm[14] ;
assign ALU_carry = \imm[15] ;
assign ALU_carry = \imm[16] ;
assign ALU_carry = \imm[17] ;
assign ALU_carry = \imm[18] ;
assign ALU_carry = \imm[19] ;
assign ALU_carry = \imm[20] ;
assign ALU_carry = \imm[21] ;
assign ALU_carry = \imm[22] ;
assign ALU_carry = \imm[23] ;
assign ALU_carry = \imm[24] ;
assign ALU_carry = \imm[25] ;
assign ALU_carry = \imm[26] ;
assign ALU_carry = \imm[27] ;
assign ALU_carry = \imm[28] ;
assign ALU_carry = \imm[29] ;
assign ALU_carry = \imm[30] ;
assign ALU_carry = \imm[31] ;
assign ALU_carry = \rd[0] ;
assign ALU_carry = \rd[1] ;
assign ALU_carry = \rd[2] ;
assign ALU_carry = \rd[3] ;
assign ALU_carry = \rd[4] ;
assign ALU_carry = \ALU_ctrl[0] ;
assign ALU_carry = \ALU_ctrl[1] ;
assign ALU_carry = \ALU_ctrl[2] ;
assign ALU_carry = \ALU_ctrl[3] ;
assign ALU_carry = \rs1_out[0] ;
assign ALU_carry = \rs1_out[1] ;
assign ALU_carry = \rs1_out[2] ;
assign ALU_carry = \rs1_out[3] ;
assign ALU_carry = \rs1_out[4] ;
assign ALU_carry = \rs1_out[5] ;
assign ALU_carry = \rs1_out[6] ;
assign ALU_carry = \rs1_out[7] ;
assign ALU_carry = \rs1_out[8] ;
assign ALU_carry = \rs1_out[9] ;
assign ALU_carry = \rs1_out[10] ;
assign ALU_carry = \rs1_out[11] ;
assign ALU_carry = \rs1_out[12] ;
assign ALU_carry = \rs1_out[13] ;
assign ALU_carry = \rs1_out[14] ;
assign ALU_carry = \rs1_out[15] ;
assign ALU_carry = \rs1_out[16] ;
assign ALU_carry = \rs1_out[17] ;
assign ALU_carry = \rs1_out[18] ;
assign ALU_carry = \rs1_out[19] ;
assign ALU_carry = \rs1_out[20] ;
assign ALU_carry = \rs1_out[21] ;
assign ALU_carry = \rs1_out[22] ;
assign ALU_carry = \rs1_out[23] ;
assign ALU_carry = \rs1_out[24] ;
assign ALU_carry = \rs1_out[25] ;
assign ALU_carry = \rs1_out[26] ;
assign ALU_carry = \rs1_out[27] ;
assign ALU_carry = \rs1_out[28] ;
assign ALU_carry = \rs1_out[29] ;
assign ALU_carry = \rs1_out[30] ;
assign ALU_carry = \rs1_out[31] ;
assign ALU_carry = \rs2_out[0] ;
assign ALU_carry = \rs2_out[1] ;
assign ALU_carry = \rs2_out[2] ;
assign ALU_carry = \rs2_out[3] ;
assign ALU_carry = \rs2_out[4] ;
assign ALU_carry = \rs2_out[5] ;
assign ALU_carry = \rs2_out[6] ;
assign ALU_carry = \rs2_out[7] ;
assign ALU_carry = \rs2_out[8] ;
assign ALU_carry = \rs2_out[9] ;
assign ALU_carry = \rs2_out[10] ;
assign ALU_carry = \rs2_out[11] ;
assign ALU_carry = \rs2_out[12] ;
assign ALU_carry = \rs2_out[13] ;
assign ALU_carry = \rs2_out[14] ;
assign ALU_carry = \rs2_out[15] ;
assign ALU_carry = \rs2_out[16] ;
assign ALU_carry = \rs2_out[17] ;
assign ALU_carry = \rs2_out[18] ;
assign ALU_carry = \rs2_out[19] ;
assign ALU_carry = \rs2_out[20] ;
assign ALU_carry = \rs2_out[21] ;
assign ALU_carry = \rs2_out[22] ;
assign ALU_carry = \rs2_out[23] ;
assign ALU_carry = \rs2_out[24] ;
assign ALU_carry = \rs2_out[25] ;
assign ALU_carry = \rs2_out[26] ;
assign ALU_carry = \rs2_out[27] ;
assign ALU_carry = \rs2_out[28] ;
assign ALU_carry = \rs2_out[29] ;
assign ALU_carry = \rs2_out[30] ;
assign ALU_carry = \rs2_out[31] ;

LOGIC0_X1 _0_ ( .Z(ALU_carry ) );

endmodule
