//Generate the verilog at 2025-08-31T15:49:25 by iSTA.
module ysyx_25030077_top (
clk,
reset,
ALU_carry,
ALU_overflow,
PC_count_o,
inst_o
);

input clk ;
input reset ;
output ALU_carry ;
output ALU_overflow ;
output [31:0] PC_count_o ;
output [31:0] inst_o ;

wire clk ;
wire reset ;
wire ALU_carry ;
wire ALU_overflow ;
wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire _167_ ;
wire _168_ ;
wire _169_ ;
wire _170_ ;
wire _171_ ;
wire _172_ ;
wire _173_ ;
wire _174_ ;
wire _175_ ;
wire _176_ ;
wire _177_ ;
wire _178_ ;
wire _179_ ;
wire _180_ ;
wire _181_ ;
wire _182_ ;
wire _183_ ;
wire _184_ ;
wire _185_ ;
wire _186_ ;
wire _187_ ;
wire _188_ ;
wire _189_ ;
wire _190_ ;
wire _191_ ;
wire _192_ ;
wire _193_ ;
wire _194_ ;
wire _195_ ;
wire _196_ ;
wire _197_ ;
wire _198_ ;
wire _199_ ;
wire _200_ ;
wire _201_ ;
wire _202_ ;
wire _203_ ;
wire _204_ ;
wire _205_ ;
wire _206_ ;
wire _207_ ;
wire _208_ ;
wire _209_ ;
wire _210_ ;
wire _211_ ;
wire _212_ ;
wire _213_ ;
wire _214_ ;
wire _215_ ;
wire _216_ ;
wire _217_ ;
wire _218_ ;
wire _219_ ;
wire _220_ ;
wire _221_ ;
wire _222_ ;
wire _223_ ;
wire _224_ ;
wire _225_ ;
wire _226_ ;
wire _227_ ;
wire _228_ ;
wire _229_ ;
wire _230_ ;
wire _231_ ;
wire _232_ ;
wire _233_ ;
wire _234_ ;
wire _235_ ;
wire _236_ ;
wire _237_ ;
wire _238_ ;
wire _239_ ;
wire _240_ ;
wire _241_ ;
wire _242_ ;
wire _243_ ;
wire _244_ ;
wire _245_ ;
wire _246_ ;
wire _247_ ;
wire _248_ ;
wire _249_ ;
wire _250_ ;
wire _251_ ;
wire _252_ ;
wire _253_ ;
wire _254_ ;
wire _255_ ;
wire _256_ ;
wire _257_ ;
wire _258_ ;
wire _259_ ;
wire _260_ ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XNOR__A_Y_$_OR__A_1_B ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_ORNOT__Y_A_$_ORNOT__Y_B_$_XOR__A_Y_$_OR__A_1_B ;
wire ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ;
wire ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ;
wire \i0.state_$_SDFFE_PP0P__Q_E ;
wire \i0.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \PC_count_o[0] ;
wire \PC_count_o[1] ;
wire \PC_count_o[2] ;
wire \PC_count_o[3] ;
wire \PC_count_o[4] ;
wire \PC_count_o[5] ;
wire \PC_count_o[6] ;
wire \PC_count_o[7] ;
wire \PC_count_o[8] ;
wire \PC_count_o[9] ;
wire \PC_count_o[10] ;
wire \PC_count_o[11] ;
wire \PC_count_o[12] ;
wire \PC_count_o[13] ;
wire \PC_count_o[14] ;
wire \PC_count_o[15] ;
wire \PC_count_o[16] ;
wire \PC_count_o[17] ;
wire \PC_count_o[18] ;
wire \PC_count_o[19] ;
wire \PC_count_o[20] ;
wire \PC_count_o[21] ;
wire \PC_count_o[22] ;
wire \PC_count_o[23] ;
wire \PC_count_o[24] ;
wire \PC_count_o[25] ;
wire \PC_count_o[26] ;
wire \PC_count_o[27] ;
wire \PC_count_o[28] ;
wire \PC_count_o[29] ;
wire \PC_count_o[30] ;
wire \PC_count_o[31] ;
wire \inst_o[0] ;
wire \inst_o[1] ;
wire \inst_o[2] ;
wire \inst_o[3] ;
wire \inst_o[4] ;
wire \inst_o[5] ;
wire \inst_o[6] ;
wire \inst_o[7] ;
wire \inst_o[8] ;
wire \inst_o[9] ;
wire \inst_o[10] ;
wire \inst_o[11] ;
wire \inst_o[12] ;
wire \inst_o[13] ;
wire \inst_o[14] ;
wire \inst_o[15] ;
wire \inst_o[16] ;
wire \inst_o[17] ;
wire \inst_o[18] ;
wire \inst_o[19] ;
wire \inst_o[20] ;
wire \inst_o[21] ;
wire \inst_o[22] ;
wire \inst_o[23] ;
wire \inst_o[24] ;
wire \inst_o[25] ;
wire \inst_o[26] ;
wire \inst_o[27] ;
wire \inst_o[28] ;
wire \inst_o[29] ;
wire \inst_o[30] ;
wire \inst_o[31] ;

assign PC_count_o[0] = \PC_count_o[0] ;
assign PC_count_o[0] = \PC_count_o[1] ;
assign PC_count_o[2] = \PC_count_o[2] ;
assign PC_count_o[3] = \PC_count_o[3] ;
assign PC_count_o[4] = \PC_count_o[4] ;
assign PC_count_o[5] = \PC_count_o[5] ;
assign PC_count_o[6] = \PC_count_o[6] ;
assign PC_count_o[7] = \PC_count_o[7] ;
assign PC_count_o[8] = \PC_count_o[8] ;
assign PC_count_o[9] = \PC_count_o[9] ;
assign PC_count_o[10] = \PC_count_o[10] ;
assign PC_count_o[11] = \PC_count_o[11] ;
assign PC_count_o[12] = \PC_count_o[12] ;
assign PC_count_o[13] = \PC_count_o[13] ;
assign PC_count_o[14] = \PC_count_o[14] ;
assign PC_count_o[15] = \PC_count_o[15] ;
assign PC_count_o[16] = \PC_count_o[16] ;
assign PC_count_o[17] = \PC_count_o[17] ;
assign PC_count_o[18] = \PC_count_o[18] ;
assign PC_count_o[19] = \PC_count_o[19] ;
assign PC_count_o[20] = \PC_count_o[20] ;
assign PC_count_o[21] = \PC_count_o[21] ;
assign PC_count_o[22] = \PC_count_o[22] ;
assign PC_count_o[23] = \PC_count_o[23] ;
assign PC_count_o[24] = \PC_count_o[24] ;
assign PC_count_o[25] = \PC_count_o[25] ;
assign PC_count_o[26] = \PC_count_o[26] ;
assign PC_count_o[27] = \PC_count_o[27] ;
assign PC_count_o[28] = \PC_count_o[28] ;
assign PC_count_o[29] = \PC_count_o[29] ;
assign PC_count_o[30] = \PC_count_o[30] ;
assign PC_count_o[31] = \PC_count_o[31] ;
assign inst_o[0] = \inst_o[0] ;
assign inst_o[0] = \inst_o[1] ;
assign inst_o[2] = \inst_o[2] ;
assign inst_o[3] = \inst_o[3] ;
assign inst_o[4] = \inst_o[4] ;
assign inst_o[5] = \inst_o[5] ;
assign inst_o[6] = \inst_o[6] ;
assign inst_o[7] = \inst_o[7] ;
assign PC_count_o[0] = \inst_o[8] ;
assign PC_count_o[0] = \inst_o[9] ;
assign PC_count_o[0] = \inst_o[10] ;
assign PC_count_o[0] = \inst_o[11] ;
assign PC_count_o[0] = \inst_o[12] ;
assign PC_count_o[0] = \inst_o[13] ;
assign PC_count_o[0] = \inst_o[14] ;
assign PC_count_o[0] = \inst_o[15] ;
assign PC_count_o[0] = \inst_o[16] ;
assign PC_count_o[0] = \inst_o[17] ;
assign PC_count_o[0] = \inst_o[18] ;
assign PC_count_o[0] = \inst_o[19] ;
assign PC_count_o[0] = \inst_o[20] ;
assign PC_count_o[0] = \inst_o[21] ;
assign PC_count_o[0] = \inst_o[22] ;
assign PC_count_o[0] = \inst_o[23] ;
assign PC_count_o[0] = \inst_o[24] ;
assign PC_count_o[0] = \inst_o[25] ;
assign PC_count_o[0] = \inst_o[26] ;
assign PC_count_o[0] = \inst_o[27] ;
assign PC_count_o[0] = \inst_o[28] ;
assign PC_count_o[0] = \inst_o[29] ;
assign PC_count_o[0] = \inst_o[30] ;
assign PC_count_o[0] = \inst_o[31] ;

AND2_X1 _261_ ( .A1(\inst_o[6] ), .A2(\inst_o[5] ), .ZN(_036_ ) );
INV_X1 _262_ ( .A(_036_ ), .ZN(_037_ ) );
NOR2_X1 _263_ ( .A1(_037_ ), .A2(\inst_o[4] ), .ZN(_038_ ) );
INV_X1 _264_ ( .A(\inst_o[2] ), .ZN(_039_ ) );
NAND2_X1 _265_ ( .A1(_039_ ), .A2(\inst_o[0] ), .ZN(_040_ ) );
NOR2_X1 _266_ ( .A1(_040_ ), .A2(\inst_o[3] ), .ZN(_041_ ) );
AND2_X2 _267_ ( .A1(_038_ ), .A2(_041_ ), .ZN(_042_ ) );
INV_X1 _268_ ( .A(_042_ ), .ZN(_043_ ) );
BUF_X2 _269_ ( .A(_043_ ), .Z(_044_ ) );
BUF_X2 _270_ ( .A(_044_ ), .Z(_045_ ) );
BUF_X2 _271_ ( .A(_038_ ), .Z(_046_ ) );
NOR2_X1 _272_ ( .A1(_039_ ), .A2(\inst_o[3] ), .ZN(_047_ ) );
AND2_X1 _273_ ( .A1(_047_ ), .A2(\inst_o[0] ), .ZN(_048_ ) );
AND2_X1 _274_ ( .A1(_046_ ), .A2(_048_ ), .ZN(_049_ ) );
NOR2_X1 _275_ ( .A1(_049_ ), .A2(reset ), .ZN(_050_ ) );
BUF_X2 _276_ ( .A(_050_ ), .Z(_051_ ) );
AND2_X4 _277_ ( .A1(\PC_count_o[3] ), .A2(\PC_count_o[2] ), .ZN(_052_ ) );
AND2_X4 _278_ ( .A1(\PC_count_o[5] ), .A2(\PC_count_o[4] ), .ZN(_053_ ) );
AND2_X4 _279_ ( .A1(_052_ ), .A2(_053_ ), .ZN(_054_ ) );
AND3_X4 _280_ ( .A1(_054_ ), .A2(\PC_count_o[7] ), .A3(\PC_count_o[6] ), .ZN(_055_ ) );
AND3_X4 _281_ ( .A1(_055_ ), .A2(\PC_count_o[9] ), .A3(\PC_count_o[8] ), .ZN(_056_ ) );
INV_X1 _282_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_057_ ) );
OAI211_X1 _283_ ( .A(_045_ ), .B(_051_ ), .C1(_056_ ), .C2(_057_ ), .ZN(_058_ ) );
AND2_X1 _284_ ( .A1(_056_ ), .A2(_057_ ), .ZN(_059_ ) );
NOR2_X1 _285_ ( .A1(_058_ ), .A2(_059_ ), .ZN(_000_ ) );
INV_X1 _286_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_060_ ) );
NAND2_X1 _287_ ( .A1(_055_ ), .A2(_060_ ), .ZN(_061_ ) );
XNOR2_X1 _288_ ( .A(_061_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_062_ ) );
NAND2_X1 _289_ ( .A1(_051_ ), .A2(_045_ ), .ZN(_063_ ) );
NOR2_X1 _290_ ( .A1(_062_ ), .A2(_063_ ), .ZN(_001_ ) );
AND3_X4 _291_ ( .A1(_056_ ), .A2(\PC_count_o[11] ), .A3(\PC_count_o[10] ), .ZN(_064_ ) );
AND3_X4 _292_ ( .A1(_064_ ), .A2(\PC_count_o[13] ), .A3(\PC_count_o[12] ), .ZN(_065_ ) );
AND3_X4 _293_ ( .A1(_065_ ), .A2(\PC_count_o[15] ), .A3(\PC_count_o[14] ), .ZN(_066_ ) );
AND2_X1 _294_ ( .A1(\PC_count_o[16] ), .A2(\PC_count_o[17] ), .ZN(_067_ ) );
AND2_X4 _295_ ( .A1(_066_ ), .A2(_067_ ), .ZN(_068_ ) );
AND2_X1 _296_ ( .A1(\PC_count_o[19] ), .A2(\PC_count_o[18] ), .ZN(_069_ ) );
AND2_X4 _297_ ( .A1(_068_ ), .A2(_069_ ), .ZN(_070_ ) );
AND2_X1 _298_ ( .A1(\PC_count_o[20] ), .A2(\PC_count_o[21] ), .ZN(_071_ ) );
AND2_X4 _299_ ( .A1(_070_ ), .A2(_071_ ), .ZN(_072_ ) );
AND2_X1 _300_ ( .A1(\PC_count_o[23] ), .A2(\PC_count_o[22] ), .ZN(_073_ ) );
AND2_X4 _301_ ( .A1(_072_ ), .A2(_073_ ), .ZN(_074_ ) );
INV_X1 _302_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_075_ ) );
AND2_X1 _303_ ( .A1(\PC_count_o[27] ), .A2(\PC_count_o[26] ), .ZN(_076_ ) );
NAND2_X1 _304_ ( .A1(\PC_count_o[24] ), .A2(\PC_count_o[25] ), .ZN(_077_ ) );
AOI21_X1 _305_ ( .A(_077_ ), .B1(_046_ ), .B2(_041_ ), .ZN(_078_ ) );
NAND4_X1 _306_ ( .A1(_074_ ), .A2(_075_ ), .A3(_076_ ), .A4(_078_ ), .ZN(_079_ ) );
INV_X16 _307_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_080_ ) );
NAND4_X1 _308_ ( .A1(_080_ ), .A2(\inst_o[7] ), .A3(\PC_count_o[14] ), .A4(\PC_count_o[11] ), .ZN(_081_ ) );
INV_X1 _309_ ( .A(\PC_count_o[15] ), .ZN(_082_ ) );
INV_X1 _310_ ( .A(\PC_count_o[13] ), .ZN(_083_ ) );
NOR3_X2 _311_ ( .A1(_081_ ), .A2(_082_ ), .A3(_083_ ), .ZN(_084_ ) );
AND3_X1 _312_ ( .A1(\PC_count_o[18] ), .A2(\PC_count_o[16] ), .A3(\PC_count_o[17] ), .ZN(_085_ ) );
AND2_X1 _313_ ( .A1(_084_ ), .A2(_085_ ), .ZN(_086_ ) );
AND3_X1 _314_ ( .A1(_086_ ), .A2(\PC_count_o[20] ), .A3(\PC_count_o[19] ), .ZN(_087_ ) );
AND3_X4 _315_ ( .A1(_087_ ), .A2(\PC_count_o[22] ), .A3(\PC_count_o[21] ), .ZN(_088_ ) );
AND2_X1 _316_ ( .A1(\PC_count_o[24] ), .A2(\PC_count_o[23] ), .ZN(_089_ ) );
AND2_X1 _317_ ( .A1(_088_ ), .A2(_089_ ), .ZN(_090_ ) );
AND3_X1 _318_ ( .A1(_090_ ), .A2(\PC_count_o[26] ), .A3(\PC_count_o[25] ), .ZN(_091_ ) );
AND2_X1 _319_ ( .A1(\PC_count_o[28] ), .A2(\PC_count_o[27] ), .ZN(_092_ ) );
AND3_X1 _320_ ( .A1(_091_ ), .A2(_042_ ), .A3(_092_ ), .ZN(_093_ ) );
INV_X1 _321_ ( .A(_093_ ), .ZN(_094_ ) );
AND3_X1 _322_ ( .A1(_079_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_094_ ), .ZN(_095_ ) );
AOI21_X1 _323_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_079_ ), .B2(_094_ ), .ZN(_096_ ) );
INV_X1 _324_ ( .A(_050_ ), .ZN(_097_ ) );
BUF_X4 _325_ ( .A(_097_ ), .Z(_098_ ) );
NOR3_X1 _326_ ( .A1(_095_ ), .A2(_096_ ), .A3(_098_ ), .ZN(_002_ ) );
AND3_X2 _327_ ( .A1(_074_ ), .A2(_076_ ), .A3(_078_ ), .ZN(_099_ ) );
INV_X1 _328_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_100_ ) );
AND3_X1 _329_ ( .A1(_091_ ), .A2(_100_ ), .A3(_042_ ), .ZN(_101_ ) );
NOR2_X1 _330_ ( .A1(_099_ ), .A2(_101_ ), .ZN(_102_ ) );
AOI21_X1 _331_ ( .A(_098_ ), .B1(_102_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_103_ ) );
OAI21_X1 _332_ ( .A(_075_ ), .B1(_099_ ), .B2(_101_ ), .ZN(_104_ ) );
AND2_X1 _333_ ( .A1(_103_ ), .A2(_104_ ), .ZN(_003_ ) );
INV_X1 _334_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_105_ ) );
NAND4_X1 _335_ ( .A1(_072_ ), .A2(_105_ ), .A3(_073_ ), .A4(_078_ ), .ZN(_106_ ) );
BUF_X4 _336_ ( .A(_042_ ), .Z(_107_ ) );
NAND4_X1 _337_ ( .A1(_090_ ), .A2(\PC_count_o[26] ), .A3(\PC_count_o[25] ), .A4(_107_ ), .ZN(_108_ ) );
NAND2_X1 _338_ ( .A1(_106_ ), .A2(_108_ ), .ZN(_109_ ) );
OAI21_X1 _339_ ( .A(_051_ ), .B1(_109_ ), .B2(_100_ ), .ZN(_110_ ) );
AND3_X1 _340_ ( .A1(_086_ ), .A2(\PC_count_o[20] ), .A3(\PC_count_o[19] ), .ZN(_111_ ) );
AND3_X1 _341_ ( .A1(_111_ ), .A2(\PC_count_o[22] ), .A3(\PC_count_o[21] ), .ZN(_112_ ) );
AND3_X1 _342_ ( .A1(_112_ ), .A2(\PC_count_o[24] ), .A3(\PC_count_o[23] ), .ZN(_113_ ) );
AND3_X1 _343_ ( .A1(_113_ ), .A2(\PC_count_o[26] ), .A3(\PC_count_o[25] ), .ZN(_114_ ) );
AND4_X1 _344_ ( .A1(_105_ ), .A2(_074_ ), .A3(\PC_count_o[24] ), .A4(\PC_count_o[25] ), .ZN(_115_ ) );
MUX2_X1 _345_ ( .A(_114_ ), .B(_115_ ), .S(_045_ ), .Z(_116_ ) );
AOI21_X1 _346_ ( .A(_110_ ), .B1(_116_ ), .B2(_100_ ), .ZN(_004_ ) );
AND2_X1 _347_ ( .A1(_074_ ), .A2(_078_ ), .ZN(_117_ ) );
INV_X1 _348_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_118_ ) );
AND4_X1 _349_ ( .A1(_118_ ), .A2(_088_ ), .A3(_042_ ), .A4(_089_ ), .ZN(_119_ ) );
OAI21_X1 _350_ ( .A(_105_ ), .B1(_117_ ), .B2(_119_ ), .ZN(_120_ ) );
AOI21_X1 _351_ ( .A(_119_ ), .B1(_074_ ), .B2(_078_ ), .ZN(_121_ ) );
AOI21_X1 _352_ ( .A(_097_ ), .B1(_121_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_122_ ) );
AND2_X1 _353_ ( .A1(_120_ ), .A2(_122_ ), .ZN(_005_ ) );
INV_X1 _354_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_123_ ) );
NAND4_X1 _355_ ( .A1(_072_ ), .A2(_123_ ), .A3(_044_ ), .A4(_073_ ), .ZN(_124_ ) );
NAND3_X1 _356_ ( .A1(_088_ ), .A2(_107_ ), .A3(_089_ ), .ZN(_125_ ) );
NAND2_X1 _357_ ( .A1(_124_ ), .A2(_125_ ), .ZN(_126_ ) );
OAI21_X1 _358_ ( .A(_051_ ), .B1(_126_ ), .B2(_118_ ), .ZN(_127_ ) );
AND4_X1 _359_ ( .A1(_123_ ), .A2(_070_ ), .A3(_073_ ), .A4(_071_ ), .ZN(_128_ ) );
MUX2_X1 _360_ ( .A(_113_ ), .B(_128_ ), .S(_045_ ), .Z(_129_ ) );
AOI21_X1 _361_ ( .A(_127_ ), .B1(_118_ ), .B2(_129_ ), .ZN(_006_ ) );
AND4_X1 _362_ ( .A1(_044_ ), .A2(_070_ ), .A3(_073_ ), .A4(_071_ ), .ZN(_130_ ) );
INV_X1 _363_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_131_ ) );
AND3_X1 _364_ ( .A1(_088_ ), .A2(_131_ ), .A3(_042_ ), .ZN(_132_ ) );
NOR2_X1 _365_ ( .A1(_130_ ), .A2(_132_ ), .ZN(_133_ ) );
AOI21_X1 _366_ ( .A(_098_ ), .B1(_133_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_134_ ) );
OAI21_X1 _367_ ( .A(_123_ ), .B1(_130_ ), .B2(_132_ ), .ZN(_135_ ) );
AND2_X1 _368_ ( .A1(_134_ ), .A2(_135_ ), .ZN(_007_ ) );
INV_X1 _369_ ( .A(_072_ ), .ZN(_136_ ) );
NOR3_X1 _370_ ( .A1(_136_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_042_ ), .ZN(_137_ ) );
AND2_X1 _371_ ( .A1(_088_ ), .A2(_042_ ), .ZN(_138_ ) );
NOR2_X1 _372_ ( .A1(_137_ ), .A2(_138_ ), .ZN(_139_ ) );
AOI21_X1 _373_ ( .A(_098_ ), .B1(_139_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_140_ ) );
AND4_X1 _374_ ( .A1(\PC_count_o[20] ), .A2(_086_ ), .A3(\PC_count_o[19] ), .A4(\PC_count_o[22] ), .ZN(_141_ ) );
AND3_X1 _375_ ( .A1(_141_ ), .A2(\PC_count_o[21] ), .A3(_042_ ), .ZN(_142_ ) );
OAI21_X1 _376_ ( .A(_131_ ), .B1(_137_ ), .B2(_142_ ), .ZN(_143_ ) );
AND2_X1 _377_ ( .A1(_140_ ), .A2(_143_ ), .ZN(_008_ ) );
NAND4_X1 _378_ ( .A1(_068_ ), .A2(_045_ ), .A3(_071_ ), .A4(_069_ ), .ZN(_144_ ) );
INV_X1 _379_ ( .A(_087_ ), .ZN(_145_ ) );
OR3_X1 _380_ ( .A1(_145_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_044_ ), .ZN(_146_ ) );
AND3_X1 _381_ ( .A1(_144_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_146_ ), .ZN(_147_ ) );
AOI21_X1 _382_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_144_ ), .B2(_146_ ), .ZN(_148_ ) );
NOR3_X1 _383_ ( .A1(_147_ ), .A2(_148_ ), .A3(_098_ ), .ZN(_009_ ) );
AOI21_X1 _384_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_046_ ), .B2(_041_ ), .ZN(_149_ ) );
NAND4_X1 _385_ ( .A1(_066_ ), .A2(_069_ ), .A3(_067_ ), .A4(_149_ ), .ZN(_150_ ) );
NAND2_X1 _386_ ( .A1(_087_ ), .A2(_107_ ), .ZN(_151_ ) );
AND3_X1 _387_ ( .A1(_150_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_151_ ), .ZN(_152_ ) );
AOI21_X1 _388_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_150_ ), .B2(_151_ ), .ZN(_153_ ) );
NOR3_X1 _389_ ( .A1(_152_ ), .A2(_153_ ), .A3(_098_ ), .ZN(_010_ ) );
AND4_X1 _390_ ( .A1(_044_ ), .A2(_066_ ), .A3(_069_ ), .A4(_067_ ), .ZN(_154_ ) );
INV_X1 _391_ ( .A(_086_ ), .ZN(_155_ ) );
NOR3_X1 _392_ ( .A1(_155_ ), .A2(_044_ ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_156_ ) );
NOR2_X1 _393_ ( .A1(_154_ ), .A2(_156_ ), .ZN(_157_ ) );
OR2_X1 _394_ ( .A1(_157_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_158_ ) );
AOI21_X1 _395_ ( .A(_097_ ), .B1(_157_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_159_ ) );
AND2_X1 _396_ ( .A1(_158_ ), .A2(_159_ ), .ZN(_011_ ) );
OAI211_X1 _397_ ( .A(_050_ ), .B(_045_ ), .C1(_060_ ), .C2(_055_ ), .ZN(_160_ ) );
AOI21_X1 _398_ ( .A(_160_ ), .B1(_060_ ), .B2(_055_ ), .ZN(_012_ ) );
INV_X1 _399_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_161_ ) );
NAND4_X1 _400_ ( .A1(_066_ ), .A2(_161_ ), .A3(_044_ ), .A4(_067_ ), .ZN(_162_ ) );
AND3_X1 _401_ ( .A1(_042_ ), .A2(_084_ ), .A3(_085_ ), .ZN(_163_ ) );
INV_X1 _402_ ( .A(_163_ ), .ZN(_164_ ) );
AND3_X1 _403_ ( .A1(_162_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_164_ ), .ZN(_165_ ) );
AOI21_X1 _404_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_162_ ), .B2(_164_ ), .ZN(_166_ ) );
NOR3_X1 _405_ ( .A1(_165_ ), .A2(_166_ ), .A3(_098_ ), .ZN(_013_ ) );
NAND3_X1 _406_ ( .A1(_066_ ), .A2(_044_ ), .A3(_067_ ), .ZN(_167_ ) );
NAND3_X1 _407_ ( .A1(_107_ ), .A2(\PC_count_o[16] ), .A3(_084_ ), .ZN(_168_ ) );
OAI21_X1 _408_ ( .A(_167_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .B2(_168_ ), .ZN(_169_ ) );
AND2_X1 _409_ ( .A1(_169_ ), .A2(_161_ ), .ZN(_170_ ) );
OAI21_X1 _410_ ( .A(_051_ ), .B1(_169_ ), .B2(_161_ ), .ZN(_171_ ) );
NOR2_X1 _411_ ( .A1(_170_ ), .A2(_171_ ), .ZN(_014_ ) );
NAND4_X1 _412_ ( .A1(_084_ ), .A2(_046_ ), .A3(\PC_count_o[16] ), .A4(_041_ ), .ZN(_172_ ) );
OAI21_X1 _413_ ( .A(_172_ ), .B1(_107_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_173_ ) );
OAI21_X1 _414_ ( .A(_173_ ), .B1(_066_ ), .B2(_107_ ), .ZN(_174_ ) );
AND2_X1 _415_ ( .A1(_174_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_175_ ) );
NOR2_X1 _416_ ( .A1(_174_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_176_ ) );
NOR3_X1 _417_ ( .A1(_175_ ), .A2(_176_ ), .A3(_098_ ), .ZN(_015_ ) );
NAND4_X1 _418_ ( .A1(_065_ ), .A2(\PC_count_o[15] ), .A3(\PC_count_o[14] ), .A4(_044_ ), .ZN(_177_ ) );
OR4_X1 _419_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(_043_ ), .A3(_083_ ), .A4(_081_ ), .ZN(_178_ ) );
NAND2_X1 _420_ ( .A1(_177_ ), .A2(_178_ ), .ZN(_179_ ) );
INV_X1 _421_ ( .A(_179_ ), .ZN(_180_ ) );
OR2_X1 _422_ ( .A1(_180_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_181_ ) );
AOI21_X1 _423_ ( .A(_097_ ), .B1(_180_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_182_ ) );
AND2_X1 _424_ ( .A1(_181_ ), .A2(_182_ ), .ZN(_016_ ) );
NOR2_X1 _425_ ( .A1(_081_ ), .A2(_083_ ), .ZN(_183_ ) );
AND3_X1 _426_ ( .A1(_046_ ), .A2(_183_ ), .A3(_041_ ), .ZN(_184_ ) );
AOI21_X1 _427_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_046_ ), .B2(_041_ ), .ZN(_185_ ) );
AOI21_X1 _428_ ( .A(_184_ ), .B1(_065_ ), .B2(_185_ ), .ZN(_186_ ) );
OAI21_X1 _429_ ( .A(_051_ ), .B1(_186_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_187_ ) );
AOI21_X1 _430_ ( .A(_187_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .B2(_186_ ), .ZN(_017_ ) );
INV_X1 _431_ ( .A(_041_ ), .ZN(_188_ ) );
AND2_X1 _432_ ( .A1(\inst_o[7] ), .A2(\PC_count_o[11] ), .ZN(_189_ ) );
AND2_X1 _433_ ( .A1(_189_ ), .A2(_080_ ), .ZN(_190_ ) );
OR4_X1 _434_ ( .A1(\inst_o[4] ), .A2(_188_ ), .A3(_037_ ), .A4(_190_ ), .ZN(_191_ ) );
NAND3_X1 _435_ ( .A1(_046_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_041_ ), .ZN(_192_ ) );
AND2_X1 _436_ ( .A1(_191_ ), .A2(_192_ ), .ZN(_193_ ) );
OAI21_X1 _437_ ( .A(_193_ ), .B1(_065_ ), .B2(_107_ ), .ZN(_194_ ) );
OAI21_X1 _438_ ( .A(_050_ ), .B1(_194_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_195_ ) );
AOI21_X1 _439_ ( .A(_195_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .B2(_194_ ), .ZN(_018_ ) );
MUX2_X1 _440_ ( .A(_189_ ), .B(_064_ ), .S(_043_ ), .Z(_196_ ) );
NOR2_X1 _441_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_197_ ) );
AND2_X1 _442_ ( .A1(_196_ ), .A2(_080_ ), .ZN(_198_ ) );
INV_X1 _443_ ( .A(_198_ ), .ZN(_199_ ) );
AOI221_X4 _444_ ( .A(_097_ ), .B1(_196_ ), .B2(_197_ ), .C1(_199_ ), .C2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_019_ ) );
OAI21_X1 _445_ ( .A(_051_ ), .B1(_196_ ), .B2(_080_ ), .ZN(_200_ ) );
NOR2_X1 _446_ ( .A1(_198_ ), .A2(_200_ ), .ZN(_020_ ) );
XNOR2_X1 _447_ ( .A(\inst_o[7] ), .B(\PC_count_o[11] ), .ZN(_201_ ) );
AND3_X1 _448_ ( .A1(_046_ ), .A2(_041_ ), .A3(_201_ ), .ZN(_202_ ) );
XOR2_X1 _449_ ( .A(_059_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .Z(_203_ ) );
AOI211_X1 _450_ ( .A(_098_ ), .B(_202_ ), .C1(_203_ ), .C2(_045_ ), .ZN(_021_ ) );
INV_X1 _451_ ( .A(_054_ ), .ZN(_204_ ) );
OR2_X1 _452_ ( .A1(_204_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_205_ ) );
XNOR2_X1 _453_ ( .A(_205_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_206_ ) );
NOR2_X1 _454_ ( .A1(_206_ ), .A2(_063_ ), .ZN(_022_ ) );
NAND2_X1 _455_ ( .A1(_204_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_207_ ) );
AND4_X1 _456_ ( .A1(_045_ ), .A2(_051_ ), .A3(_205_ ), .A4(_207_ ), .ZN(_023_ ) );
INV_X1 _457_ ( .A(_052_ ), .ZN(_208_ ) );
OAI21_X1 _458_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .B1(_208_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_209_ ) );
OR3_X1 _459_ ( .A1(_208_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_210_ ) );
AND4_X1 _460_ ( .A1(_045_ ), .A2(_051_ ), .A3(_209_ ), .A4(_210_ ), .ZN(_024_ ) );
XOR2_X1 _461_ ( .A(_052_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .Z(_211_ ) );
NOR4_X1 _462_ ( .A1(_107_ ), .A2(_049_ ), .A3(_211_ ), .A4(reset ), .ZN(_025_ ) );
INV_X1 _463_ ( .A(\PC_count_o[3] ), .ZN(_212_ ) );
INV_X1 _464_ ( .A(\PC_count_o[2] ), .ZN(_213_ ) );
NAND2_X1 _465_ ( .A1(_212_ ), .A2(_213_ ), .ZN(_214_ ) );
AND4_X1 _466_ ( .A1(_208_ ), .A2(_051_ ), .A3(_045_ ), .A4(_214_ ), .ZN(_026_ ) );
NOR4_X1 _467_ ( .A1(_107_ ), .A2(_049_ ), .A3(reset ), .A4(\PC_count_o[2] ), .ZN(_027_ ) );
AND3_X1 _468_ ( .A1(_076_ ), .A2(\PC_count_o[29] ), .A3(\PC_count_o[28] ), .ZN(_215_ ) );
AND3_X4 _469_ ( .A1(_074_ ), .A2(_078_ ), .A3(_215_ ), .ZN(_216_ ) );
INV_X1 _470_ ( .A(_091_ ), .ZN(_217_ ) );
INV_X1 _471_ ( .A(_092_ ), .ZN(_218_ ) );
NOR4_X1 _472_ ( .A1(_217_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_044_ ), .A4(_218_ ), .ZN(_219_ ) );
NOR2_X1 _473_ ( .A1(_216_ ), .A2(_219_ ), .ZN(_220_ ) );
AOI21_X1 _474_ ( .A(_098_ ), .B1(_220_ ), .B2(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_221_ ) );
INV_X1 _475_ ( .A(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_222_ ) );
OAI21_X1 _476_ ( .A(_222_ ), .B1(_216_ ), .B2(_219_ ), .ZN(_223_ ) );
AND2_X1 _477_ ( .A1(_221_ ), .A2(_223_ ), .ZN(_028_ ) );
INV_X1 _478_ ( .A(reset ), .ZN(_224_ ) );
NAND4_X4 _479_ ( .A1(_074_ ), .A2(_222_ ), .A3(_078_ ), .A4(_215_ ), .ZN(_225_ ) );
NAND3_X1 _480_ ( .A1(_093_ ), .A2(\PC_count_o[29] ), .A3(\PC_count_o[30] ), .ZN(_226_ ) );
AND2_X2 _481_ ( .A1(_225_ ), .A2(_226_ ), .ZN(_227_ ) );
XNOR2_X2 _482_ ( .A(_227_ ), .B(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_228_ ) );
OAI21_X1 _483_ ( .A(_224_ ), .B1(_228_ ), .B2(_049_ ), .ZN(_029_ ) );
AND2_X1 _484_ ( .A1(_224_ ), .A2(\PC_count_o[7] ), .ZN(_030_ ) );
AND2_X1 _485_ ( .A1(_224_ ), .A2(\PC_count_o[6] ), .ZN(_031_ ) );
AND2_X1 _486_ ( .A1(_224_ ), .A2(\PC_count_o[5] ), .ZN(_032_ ) );
AND2_X1 _487_ ( .A1(_224_ ), .A2(\PC_count_o[4] ), .ZN(_033_ ) );
NOR2_X1 _488_ ( .A1(_212_ ), .A2(reset ), .ZN(_034_ ) );
NOR2_X1 _489_ ( .A1(_213_ ), .A2(reset ), .ZN(_035_ ) );
XOR2_X1 _490_ ( .A(\inst_o[5] ), .B(\inst_o[4] ), .Z(_229_ ) );
OR3_X1 _491_ ( .A1(_188_ ), .A2(_229_ ), .A3(\inst_o[6] ), .ZN(_230_ ) );
OR4_X1 _492_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_231_ ) );
NOR4_X1 _493_ ( .A1(_231_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_232_ ) );
NOR4_X1 _494_ ( .A1(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_233_ ) );
NOR4_X1 _495_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_234_ ) );
AND3_X1 _496_ ( .A1(_232_ ), .A2(_233_ ), .A3(_234_ ), .ZN(_235_ ) );
AND2_X1 _497_ ( .A1(\inst_o[2] ), .A2(\inst_o[0] ), .ZN(_236_ ) );
AND2_X1 _498_ ( .A1(_046_ ), .A2(_236_ ), .ZN(_237_ ) );
INV_X1 _499_ ( .A(_237_ ), .ZN(_238_ ) );
NOR2_X1 _500_ ( .A1(\inst_o[6] ), .A2(\inst_o[5] ), .ZN(_239_ ) );
NAND3_X1 _501_ ( .A1(_048_ ), .A2(\inst_o[4] ), .A3(_239_ ), .ZN(_240_ ) );
AOI21_X1 _502_ ( .A(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_238_ ), .B2(_240_ ), .ZN(_241_ ) );
NOR4_X1 _503_ ( .A1(_082_ ), .A2(_212_ ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ), .ZN(_242_ ) );
NOR4_X1 _504_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_243_ ) );
NOR4_X1 _505_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_244_ ) );
AND4_X1 _506_ ( .A1(_197_ ), .A2(_242_ ), .A3(_243_ ), .A4(_244_ ), .ZN(_245_ ) );
AND2_X1 _507_ ( .A1(_245_ ), .A2(_237_ ), .ZN(_246_ ) );
AND4_X1 _508_ ( .A1(_230_ ), .A2(_235_ ), .A3(_241_ ), .A4(_246_ ), .ZN(ALU_carry ) );
INV_X1 _509_ ( .A(_246_ ), .ZN(_247_ ) );
NAND4_X1 _510_ ( .A1(_230_ ), .A2(_232_ ), .A3(_233_ ), .A4(_234_ ), .ZN(_248_ ) );
NOR3_X1 _511_ ( .A1(_247_ ), .A2(_241_ ), .A3(_248_ ), .ZN(ALU_overflow ) );
AND3_X1 _512_ ( .A1(_046_ ), .A2(\inst_o[3] ), .A3(_236_ ), .ZN(_249_ ) );
INV_X1 _513_ ( .A(\inst_o[7] ), .ZN(_250_ ) );
NAND4_X1 _514_ ( .A1(_250_ ), .A2(\inst_o[6] ), .A3(\inst_o[5] ), .A4(\inst_o[4] ), .ZN(_251_ ) );
NOR3_X1 _515_ ( .A1(_251_ ), .A2(_040_ ), .A3(\inst_o[3] ), .ZN(_252_ ) );
NOR3_X1 _516_ ( .A1(_249_ ), .A2(_107_ ), .A3(_252_ ), .ZN(\i0.state_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _517_ ( .A1(_249_ ), .A2(_252_ ), .ZN(\i0.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
CLKGATE_X1 _518_ ( .CK(clk ), .E(\i0.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_253_ ) );
CLKGATE_X1 _519_ ( .CK(clk ), .E(\i0.state_$_SDFFE_PP0P__Q_E ), .GCK(_254_ ) );
LOGIC0_X1 _520_ ( .Z(\PC_count_o[0] ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q ( .D(_000_ ), .CK(_254_ ), .Q(\PC_count_o[10] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_1 ( .D(_001_ ), .CK(_254_ ), .Q(\PC_count_o[9] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_10 ( .D(_002_ ), .CK(_253_ ), .Q(\PC_count_o[29] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_11 ( .D(_003_ ), .CK(_253_ ), .Q(\PC_count_o[28] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_12 ( .D(_004_ ), .CK(_253_ ), .Q(\PC_count_o[27] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_13 ( .D(_005_ ), .CK(_253_ ), .Q(\PC_count_o[26] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_14 ( .D(_006_ ), .CK(_253_ ), .Q(\PC_count_o[25] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_15 ( .D(_007_ ), .CK(_253_ ), .Q(\PC_count_o[24] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_16 ( .D(_008_ ), .CK(_253_ ), .Q(\PC_count_o[23] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_17 ( .D(_009_ ), .CK(_253_ ), .Q(\PC_count_o[22] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_18 ( .D(_010_ ), .CK(_253_ ), .Q(\PC_count_o[21] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_19 ( .D(_011_ ), .CK(_253_ ), .Q(\PC_count_o[20] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_2 ( .D(_012_ ), .CK(_254_ ), .Q(\PC_count_o[8] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_20 ( .D(_013_ ), .CK(_253_ ), .Q(\PC_count_o[19] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_21 ( .D(_014_ ), .CK(_253_ ), .Q(\PC_count_o[18] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_22 ( .D(_015_ ), .CK(_253_ ), .Q(\PC_count_o[17] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_23 ( .D(_016_ ), .CK(_253_ ), .Q(\PC_count_o[16] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_24 ( .D(_017_ ), .CK(_253_ ), .Q(\PC_count_o[15] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_25 ( .D(_018_ ), .CK(_253_ ), .Q(\PC_count_o[14] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_26 ( .D(_019_ ), .CK(_253_ ), .Q(\PC_count_o[13] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_27 ( .D(_020_ ), .CK(_253_ ), .Q(\PC_count_o[12] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_28 ( .D(_021_ ), .CK(_253_ ), .Q(\PC_count_o[11] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_3 ( .D(_022_ ), .CK(_254_ ), .Q(\PC_count_o[7] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_4 ( .D(_023_ ), .CK(_254_ ), .Q(\PC_count_o[6] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_5 ( .D(_024_ ), .CK(_254_ ), .Q(\PC_count_o[5] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_6 ( .D(_025_ ), .CK(_254_ ), .Q(\PC_count_o[4] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_7 ( .D(_026_ ), .CK(_254_ ), .Q(\PC_count_o[3] ), .QN(_260_ ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_8 ( .D(_027_ ), .CK(_254_ ), .Q(\PC_count_o[2] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_9 ( .D(_028_ ), .CK(_253_ ), .Q(\PC_count_o[30] ), .QN(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP1P__Q ( .D(_029_ ), .CK(_253_ ), .Q(\PC_count_o[31] ), .QN(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q ( .D(_030_ ), .CK(clk ), .Q(\inst_o[7] ), .QN(_259_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_1 ( .D(_031_ ), .CK(clk ), .Q(\inst_o[6] ), .QN(_258_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_2 ( .D(_032_ ), .CK(clk ), .Q(\inst_o[5] ), .QN(_257_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_3 ( .D(_033_ ), .CK(clk ), .Q(\inst_o[4] ), .QN(_256_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_4 ( .D(_034_ ), .CK(clk ), .Q(\inst_o[3] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XNOR__A_Y_$_OR__A_1_B ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_5 ( .D(_035_ ), .CK(clk ), .Q(\inst_o[2] ), .QN(_255_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_6 ( .D(\PC_count_o[0] ), .CK(clk ), .Q(\inst_o[0] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_ORNOT__Y_A_$_ORNOT__Y_B_$_XOR__A_Y_$_OR__A_1_B ) );

endmodule
