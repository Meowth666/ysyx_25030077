//Generate the verilog at 2025-09-25T17:34:57 by iSTA.
module top (
clock,
reset,
io_is_unknown_instruction,
io_carry,
io_isoverflow
);

input clock ;
input reset ;
output io_is_unknown_instruction ;
output io_carry ;
output io_isoverflow ;

wire clock ;
wire reset ;
wire io_is_unknown_instruction ;
wire io_carry ;
wire io_isoverflow ;
wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire \b_ifu.io_ar_ready ;
wire \b_ifu.io_ar_valid ;
wire \b_ifu.io_rd_Req_valid ;
wire \b_ifu.reqQ.maybe_full_$_SDFFE_PP0P__Q_E ;
wire \c_arbiter._inst_reg_T_2 ;
wire \c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ;
wire \c_arbiter.io_axi_b_ready ;
wire \f_gpr.canAccept_prng.state_0_$_DFF_P__Q_D ;
wire \g_mem._startDelay_T ;
wire \g_mem.canAccept_prng.state_0_$_DFF_P__Q_D ;
wire \g_mem.delayCnt_prng.state_0_$_DFF_P__Q_D ;
wire \g_mem.validReg ;
wire [2:0] \c_arbiter.inst_reg ;
wire [2:0] \c_arbiter.io_axi_r_data ;
wire [2:0] \c_arbiter.io_delay_cnt ;
wire [1:0] \c_arbiter.state_reg ;
wire [15:0] \f_gpr._canAccept_T ;
wire [15:0] \g_mem._canAccept_T ;
wire [2:0] \g_mem._delayCnt_T ;

assign io_isoverflow = io_carry ;

INV_X1 _147_ ( .A(\b_ifu.io_rd_Req_valid ), .ZN(_046_ ) );
NOR3_X1 _148_ ( .A1(_046_ ), .A2(reset ), .A3(\b_ifu.io_ar_valid ), .ZN(_000_ ) );
INV_X1 _149_ ( .A(reset ), .ZN(_047_ ) );
CLKBUF_X2 _150_ ( .A(_047_ ), .Z(_044_ ) );
AND2_X1 _151_ ( .A1(_044_ ), .A2(\c_arbiter.io_axi_r_data [2] ), .ZN(_001_ ) );
AND2_X1 _152_ ( .A1(_044_ ), .A2(\c_arbiter.io_axi_r_data [1] ), .ZN(_002_ ) );
AND2_X1 _153_ ( .A1(_044_ ), .A2(\c_arbiter.io_axi_r_data [0] ), .ZN(_003_ ) );
NAND2_X4 _154_ ( .A1(\c_arbiter.inst_reg [0] ), .A2(\c_arbiter.inst_reg [1] ), .ZN(_048_ ) );
OR2_X2 _155_ ( .A1(_048_ ), .A2(\c_arbiter.inst_reg [2] ), .ZN(io_is_unknown_instruction ) );
AOI211_X1 _156_ ( .A(reset ), .B(\c_arbiter.state_reg [1] ), .C1(io_is_unknown_instruction ), .C2(\c_arbiter.state_reg [0] ), .ZN(_004_ ) );
NOR2_X4 _157_ ( .A1(\c_arbiter.io_delay_cnt [1] ), .A2(\c_arbiter.io_delay_cnt [0] ), .ZN(_049_ ) );
AND2_X4 _158_ ( .A1(_049_ ), .A2(\c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ), .ZN(_050_ ) );
NAND4_X1 _159_ ( .A1(_050_ ), .A2(io_is_unknown_instruction ), .A3(\b_ifu.io_ar_ready ), .A4(\g_mem.validReg ), .ZN(_051_ ) );
INV_X16 _160_ ( .A(\c_arbiter.state_reg [1] ), .ZN(_052_ ) );
AND2_X4 _161_ ( .A1(_052_ ), .A2(\c_arbiter.state_reg [0] ), .ZN(_053_ ) );
INV_X1 _162_ ( .A(\c_arbiter.io_delay_cnt [1] ), .ZN(_054_ ) );
AND3_X1 _163_ ( .A1(_054_ ), .A2(\c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ), .A3(\c_arbiter.io_delay_cnt [0] ), .ZN(_055_ ) );
INV_X1 _164_ ( .A(_055_ ), .ZN(_056_ ) );
OAI211_X1 _165_ ( .A(_051_ ), .B(_053_ ), .C1(io_is_unknown_instruction ), .C2(_056_ ), .ZN(_057_ ) );
NOR2_X1 _166_ ( .A1(\c_arbiter.state_reg [1] ), .A2(\c_arbiter.state_reg [0] ), .ZN(_058_ ) );
AND4_X1 _167_ ( .A1(\c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ), .A2(_058_ ), .A3(_054_ ), .A4(\c_arbiter.io_delay_cnt [0] ), .ZN(\c_arbiter._inst_reg_T_2 ) );
INV_X1 _168_ ( .A(\c_arbiter._inst_reg_T_2 ), .ZN(_059_ ) );
AOI21_X1 _169_ ( .A(reset ), .B1(_057_ ), .B2(_059_ ), .ZN(_005_ ) );
AND2_X1 _170_ ( .A1(_050_ ), .A2(\g_mem.validReg ), .ZN(_060_ ) );
AND2_X1 _171_ ( .A1(_060_ ), .A2(\b_ifu.io_ar_ready ), .ZN(_061_ ) );
OR3_X1 _172_ ( .A1(_061_ ), .A2(_052_ ), .A3(\c_arbiter.state_reg [0] ), .ZN(_062_ ) );
OAI21_X1 _173_ ( .A(_051_ ), .B1(io_is_unknown_instruction ), .B2(_056_ ), .ZN(_063_ ) );
NAND2_X1 _174_ ( .A1(_063_ ), .A2(_053_ ), .ZN(_064_ ) );
AOI21_X1 _175_ ( .A(reset ), .B1(_062_ ), .B2(_064_ ), .ZN(_006_ ) );
AND2_X1 _176_ ( .A1(_044_ ), .A2(\f_gpr._canAccept_T [9] ), .ZN(_007_ ) );
AND2_X1 _177_ ( .A1(_044_ ), .A2(\f_gpr._canAccept_T [10] ), .ZN(_008_ ) );
AND2_X1 _178_ ( .A1(_044_ ), .A2(\f_gpr._canAccept_T [11] ), .ZN(_009_ ) );
AND2_X1 _179_ ( .A1(_044_ ), .A2(\f_gpr._canAccept_T [12] ), .ZN(_010_ ) );
CLKBUF_X2 _180_ ( .A(_047_ ), .Z(_065_ ) );
AND2_X1 _181_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [13] ), .ZN(_011_ ) );
AND2_X1 _182_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [14] ), .ZN(_012_ ) );
INV_X1 _183_ ( .A(\c_arbiter.io_axi_b_ready ), .ZN(_066_ ) );
NOR2_X1 _184_ ( .A1(_066_ ), .A2(reset ), .ZN(_013_ ) );
AND2_X1 _185_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [1] ), .ZN(_014_ ) );
AND2_X1 _186_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [2] ), .ZN(_015_ ) );
AND2_X1 _187_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [3] ), .ZN(_016_ ) );
AND2_X1 _188_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [4] ), .ZN(_017_ ) );
AND2_X1 _189_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [5] ), .ZN(_018_ ) );
AND2_X1 _190_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [6] ), .ZN(_019_ ) );
AND2_X1 _191_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [7] ), .ZN(_020_ ) );
AND2_X1 _192_ ( .A1(_065_ ), .A2(\f_gpr._canAccept_T [8] ), .ZN(_021_ ) );
NOR3_X1 _193_ ( .A1(_066_ ), .A2(_052_ ), .A3(\c_arbiter.state_reg [0] ), .ZN(_067_ ) );
NAND3_X1 _194_ ( .A1(_050_ ), .A2(\g_mem.validReg ), .A3(_067_ ), .ZN(_068_ ) );
INV_X1 _195_ ( .A(\b_ifu.io_ar_valid ), .ZN(_069_ ) );
OAI211_X1 _196_ ( .A(_068_ ), .B(_044_ ), .C1(_046_ ), .C2(_069_ ), .ZN(_022_ ) );
CLKBUF_X2 _197_ ( .A(_047_ ), .Z(_070_ ) );
AND2_X1 _198_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [9] ), .ZN(_023_ ) );
AND2_X1 _199_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [10] ), .ZN(_024_ ) );
AND2_X1 _200_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [11] ), .ZN(_025_ ) );
AND2_X1 _201_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [12] ), .ZN(_026_ ) );
AND2_X1 _202_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [13] ), .ZN(_027_ ) );
AND2_X1 _203_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [14] ), .ZN(_028_ ) );
AND2_X1 _204_ ( .A1(_070_ ), .A2(\b_ifu.io_ar_ready ), .ZN(_029_ ) );
AND2_X1 _205_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [1] ), .ZN(_030_ ) );
AND2_X1 _206_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [2] ), .ZN(_031_ ) );
AND2_X1 _207_ ( .A1(_070_ ), .A2(\g_mem._canAccept_T [3] ), .ZN(_032_ ) );
AND2_X1 _208_ ( .A1(_047_ ), .A2(\g_mem._canAccept_T [4] ), .ZN(_033_ ) );
AND2_X1 _209_ ( .A1(_047_ ), .A2(\g_mem._canAccept_T [5] ), .ZN(_034_ ) );
AND2_X1 _210_ ( .A1(_047_ ), .A2(\g_mem._canAccept_T [6] ), .ZN(_035_ ) );
AND2_X1 _211_ ( .A1(_047_ ), .A2(\g_mem._canAccept_T [7] ), .ZN(_036_ ) );
AND2_X1 _212_ ( .A1(_047_ ), .A2(\g_mem._canAccept_T [8] ), .ZN(_037_ ) );
NAND4_X4 _213_ ( .A1(_053_ ), .A2(\c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ), .A3(\g_mem.validReg ), .A4(_049_ ), .ZN(_071_ ) );
NAND2_X1 _214_ ( .A1(_058_ ), .A2(\b_ifu.io_ar_valid ), .ZN(_072_ ) );
NAND2_X4 _215_ ( .A1(_071_ ), .A2(_072_ ), .ZN(_073_ ) );
NAND2_X4 _216_ ( .A1(_073_ ), .A2(\b_ifu.io_ar_ready ), .ZN(_074_ ) );
INV_X4 _217_ ( .A(_074_ ), .ZN(\g_mem._startDelay_T ) );
AOI21_X4 _218_ ( .A(\c_arbiter.state_reg [1] ), .B1(io_is_unknown_instruction ), .B2(\c_arbiter.state_reg [0] ), .ZN(_075_ ) );
AND2_X2 _219_ ( .A1(\g_mem._startDelay_T ), .A2(_075_ ), .ZN(_076_ ) );
INV_X1 _220_ ( .A(\c_arbiter.io_delay_cnt [0] ), .ZN(_077_ ) );
OAI211_X1 _221_ ( .A(_054_ ), .B(_077_ ), .C1(\c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ), .C2(\c_arbiter.io_delay_cnt [2] ), .ZN(_078_ ) );
OAI21_X1 _222_ ( .A(_078_ ), .B1(\c_arbiter.io_delay_cnt [2] ), .B2(_049_ ), .ZN(_079_ ) );
OR2_X2 _223_ ( .A1(_076_ ), .A2(_079_ ), .ZN(_080_ ) );
NAND4_X1 _224_ ( .A1(_073_ ), .A2(\b_ifu.io_ar_ready ), .A3(\g_mem._delayCnt_T [2] ), .A4(_075_ ), .ZN(_081_ ) );
AOI21_X1 _225_ ( .A(reset ), .B1(_080_ ), .B2(_081_ ), .ZN(_038_ ) );
AND3_X1 _226_ ( .A1(_054_ ), .A2(_077_ ), .A3(\c_arbiter.io_delay_cnt [2] ), .ZN(_082_ ) );
AOI221_X2 _227_ ( .A(_082_ ), .B1(\c_arbiter.io_delay_cnt [1] ), .B2(\c_arbiter.io_delay_cnt [0] ), .C1(\g_mem._startDelay_T ), .C2(_075_ ), .ZN(_083_ ) );
INV_X1 _228_ ( .A(\g_mem._delayCnt_T [1] ), .ZN(_084_ ) );
AOI211_X1 _229_ ( .A(reset ), .B(_083_ ), .C1(_084_ ), .C2(_076_ ), .ZN(_039_ ) );
INV_X1 _230_ ( .A(_050_ ), .ZN(_085_ ) );
AOI22_X1 _231_ ( .A1(\g_mem._startDelay_T ), .A2(_075_ ), .B1(_077_ ), .B2(_085_ ), .ZN(_086_ ) );
INV_X1 _232_ ( .A(\g_mem._delayCnt_T [0] ), .ZN(_087_ ) );
AOI211_X1 _233_ ( .A(reset ), .B(_086_ ), .C1(_087_ ), .C2(_076_ ), .ZN(_040_ ) );
NOR2_X1 _234_ ( .A1(_087_ ), .A2(reset ), .ZN(_041_ ) );
NOR2_X1 _235_ ( .A1(_084_ ), .A2(reset ), .ZN(_042_ ) );
NOR3_X1 _236_ ( .A1(reset ), .A2(\c_arbiter.state_reg [1] ), .A3(\c_arbiter.state_reg [0] ), .ZN(_043_ ) );
OAI21_X1 _237_ ( .A(\g_mem.validReg ), .B1(_085_ ), .B2(_066_ ), .ZN(_088_ ) );
AOI21_X1 _238_ ( .A(reset ), .B1(_074_ ), .B2(_088_ ), .ZN(_045_ ) );
XOR2_X1 _239_ ( .A(\f_gpr._canAccept_T [10] ), .B(\f_gpr._canAccept_T [12] ), .Z(_089_ ) );
XNOR2_X1 _240_ ( .A(\f_gpr._canAccept_T [13] ), .B(\f_gpr._canAccept_T [15] ), .ZN(_090_ ) );
AOI21_X1 _241_ ( .A(reset ), .B1(_089_ ), .B2(_090_ ), .ZN(_091_ ) );
OAI21_X1 _242_ ( .A(_091_ ), .B1(_090_ ), .B2(_089_ ), .ZN(\f_gpr.canAccept_prng.state_0_$_DFF_P__Q_D ) );
MUX2_X1 _243_ ( .A(\b_ifu.io_rd_Req_valid ), .B(\b_ifu.io_ar_ready ), .S(\b_ifu.io_ar_valid ), .Z(\b_ifu.reqQ.maybe_full_$_SDFFE_PP0P__Q_E ) );
XOR2_X1 _244_ ( .A(\g_mem._canAccept_T [10] ), .B(\g_mem._canAccept_T [12] ), .Z(_092_ ) );
XNOR2_X1 _245_ ( .A(\g_mem._canAccept_T [13] ), .B(\g_mem._canAccept_T [15] ), .ZN(_093_ ) );
AOI21_X1 _246_ ( .A(reset ), .B1(_092_ ), .B2(_093_ ), .ZN(_094_ ) );
OAI21_X1 _247_ ( .A(_094_ ), .B1(_093_ ), .B2(_092_ ), .ZN(\g_mem.canAccept_prng.state_0_$_DFF_P__Q_D ) );
XNOR2_X1 _248_ ( .A(\g_mem._delayCnt_T [1] ), .B(\g_mem._delayCnt_T [2] ), .ZN(_095_ ) );
NAND2_X1 _249_ ( .A1(_095_ ), .A2(_044_ ), .ZN(\g_mem.delayCnt_prng.state_0_$_DFF_P__Q_D ) );
CLKGATE_X1 _250_ ( .CK(clock ), .E(\g_mem._startDelay_T ), .GCK(_096_ ) );
CLKGATE_X1 _251_ ( .CK(clock ), .E(\c_arbiter._inst_reg_T_2 ), .GCK(_097_ ) );
CLKGATE_X1 _252_ ( .CK(clock ), .E(\b_ifu.reqQ.maybe_full_$_SDFFE_PP0P__Q_E ), .GCK(_098_ ) );
LOGIC0_X1 _253_ ( .Z(io_carry ) );
DFF_X1 \b_ifu.reqQ.maybe_full_$_SDFFE_PP0P__Q ( .D(_000_ ), .CK(_098_ ), .Q(\b_ifu.io_ar_valid ), .QN(_143_ ) );
DFF_X1 \c_arbiter.inst_reg_$_SDFFE_PP0P__Q ( .D(_001_ ), .CK(_097_ ), .Q(\c_arbiter.inst_reg [2] ), .QN(_142_ ) );
DFF_X1 \c_arbiter.inst_reg_$_SDFFE_PP0P__Q_1 ( .D(_002_ ), .CK(_097_ ), .Q(\c_arbiter.inst_reg [1] ), .QN(_141_ ) );
DFF_X1 \c_arbiter.inst_reg_$_SDFFE_PP0P__Q_2 ( .D(_003_ ), .CK(_097_ ), .Q(\c_arbiter.inst_reg [0] ), .QN(_140_ ) );
DFF_X1 \c_arbiter.state_reg_$_SDFF_PP0__Q ( .D(_005_ ), .CK(clock ), .Q(\c_arbiter.state_reg [0] ), .QN(_138_ ) );
DFF_X1 \c_arbiter.state_reg_$_SDFF_PP0__Q_1 ( .D(_006_ ), .CK(clock ), .Q(\c_arbiter.state_reg [1] ), .QN(_144_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_0_$_DFF_P__Q ( .D(\f_gpr.canAccept_prng.state_0_$_DFF_P__Q_D ), .CK(clock ), .Q(\c_arbiter.io_axi_b_ready ), .QN(_137_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_10_$_SDFF_PP0__Q ( .D(_007_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [10] ), .QN(_136_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_11_$_SDFF_PP0__Q ( .D(_008_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [11] ), .QN(_135_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_12_$_SDFF_PP0__Q ( .D(_009_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [12] ), .QN(_134_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_13_$_SDFF_PP0__Q ( .D(_010_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [13] ), .QN(_133_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_14_$_SDFF_PP0__Q ( .D(_011_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [14] ), .QN(_132_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_15_$_SDFF_PP0__Q ( .D(_012_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [15] ), .QN(_131_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_1_$_SDFF_PP0__Q ( .D(_013_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [1] ), .QN(_130_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_2_$_SDFF_PP0__Q ( .D(_014_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [2] ), .QN(_129_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_3_$_SDFF_PP0__Q ( .D(_015_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [3] ), .QN(_128_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_4_$_SDFF_PP0__Q ( .D(_016_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [4] ), .QN(_127_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_5_$_SDFF_PP0__Q ( .D(_017_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [5] ), .QN(_126_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_6_$_SDFF_PP0__Q ( .D(_018_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [6] ), .QN(_125_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_7_$_SDFF_PP0__Q ( .D(_019_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [7] ), .QN(_124_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_8_$_SDFF_PP0__Q ( .D(_020_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [8] ), .QN(_123_ ) );
DFF_X1 \f_gpr.canAccept_prng.state_9_$_SDFF_PP0__Q ( .D(_021_ ), .CK(clock ), .Q(\f_gpr._canAccept_T [9] ), .QN(_122_ ) );
DFF_X1 \f_gpr.validReg_$_SDFF_PP1__Q ( .D(_022_ ), .CK(clock ), .Q(\b_ifu.io_rd_Req_valid ), .QN(_145_ ) );
DFF_X1 \g_mem.canAccept_prng.state_0_$_DFF_P__Q ( .D(\g_mem.canAccept_prng.state_0_$_DFF_P__Q_D ), .CK(clock ), .Q(\b_ifu.io_ar_ready ), .QN(_121_ ) );
DFF_X1 \g_mem.canAccept_prng.state_10_$_SDFF_PP0__Q ( .D(_023_ ), .CK(clock ), .Q(\g_mem._canAccept_T [10] ), .QN(_120_ ) );
DFF_X1 \g_mem.canAccept_prng.state_11_$_SDFF_PP0__Q ( .D(_024_ ), .CK(clock ), .Q(\g_mem._canAccept_T [11] ), .QN(_119_ ) );
DFF_X1 \g_mem.canAccept_prng.state_12_$_SDFF_PP0__Q ( .D(_025_ ), .CK(clock ), .Q(\g_mem._canAccept_T [12] ), .QN(_118_ ) );
DFF_X1 \g_mem.canAccept_prng.state_13_$_SDFF_PP0__Q ( .D(_026_ ), .CK(clock ), .Q(\g_mem._canAccept_T [13] ), .QN(_117_ ) );
DFF_X1 \g_mem.canAccept_prng.state_14_$_SDFF_PP0__Q ( .D(_027_ ), .CK(clock ), .Q(\g_mem._canAccept_T [14] ), .QN(_116_ ) );
DFF_X1 \g_mem.canAccept_prng.state_15_$_SDFF_PP0__Q ( .D(_028_ ), .CK(clock ), .Q(\g_mem._canAccept_T [15] ), .QN(_115_ ) );
DFF_X1 \g_mem.canAccept_prng.state_1_$_SDFF_PP0__Q ( .D(_029_ ), .CK(clock ), .Q(\g_mem._canAccept_T [1] ), .QN(_114_ ) );
DFF_X1 \g_mem.canAccept_prng.state_2_$_SDFF_PP0__Q ( .D(_030_ ), .CK(clock ), .Q(\g_mem._canAccept_T [2] ), .QN(_113_ ) );
DFF_X1 \g_mem.canAccept_prng.state_3_$_SDFF_PP0__Q ( .D(_031_ ), .CK(clock ), .Q(\g_mem._canAccept_T [3] ), .QN(_112_ ) );
DFF_X1 \g_mem.canAccept_prng.state_4_$_SDFF_PP0__Q ( .D(_032_ ), .CK(clock ), .Q(\g_mem._canAccept_T [4] ), .QN(_111_ ) );
DFF_X1 \g_mem.canAccept_prng.state_5_$_SDFF_PP0__Q ( .D(_033_ ), .CK(clock ), .Q(\g_mem._canAccept_T [5] ), .QN(_110_ ) );
DFF_X1 \g_mem.canAccept_prng.state_6_$_SDFF_PP0__Q ( .D(_034_ ), .CK(clock ), .Q(\g_mem._canAccept_T [6] ), .QN(_109_ ) );
DFF_X1 \g_mem.canAccept_prng.state_7_$_SDFF_PP0__Q ( .D(_035_ ), .CK(clock ), .Q(\g_mem._canAccept_T [7] ), .QN(_108_ ) );
DFF_X1 \g_mem.canAccept_prng.state_8_$_SDFF_PP0__Q ( .D(_036_ ), .CK(clock ), .Q(\g_mem._canAccept_T [8] ), .QN(_107_ ) );
DFF_X1 \g_mem.canAccept_prng.state_9_$_SDFF_PP0__Q ( .D(_037_ ), .CK(clock ), .Q(\g_mem._canAccept_T [9] ), .QN(_106_ ) );
DFF_X1 \g_mem.delayCnt_$_SDFF_PP0__Q ( .D(_038_ ), .CK(clock ), .Q(\c_arbiter.io_delay_cnt [2] ), .QN(\c_arbiter._inst_reg_T_2_$_AND__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \g_mem.delayCnt_$_SDFF_PP0__Q_1 ( .D(_039_ ), .CK(clock ), .Q(\c_arbiter.io_delay_cnt [1] ), .QN(_105_ ) );
DFF_X1 \g_mem.delayCnt_$_SDFF_PP0__Q_2 ( .D(_040_ ), .CK(clock ), .Q(\c_arbiter.io_delay_cnt [0] ), .QN(_146_ ) );
DFF_X1 \g_mem.delayCnt_prng.state_0_$_DFF_P__Q ( .D(\g_mem.delayCnt_prng.state_0_$_DFF_P__Q_D ), .CK(clock ), .Q(\g_mem._delayCnt_T [0] ), .QN(_104_ ) );
DFF_X1 \g_mem.delayCnt_prng.state_1_$_SDFF_PP0__Q ( .D(_041_ ), .CK(clock ), .Q(\g_mem._delayCnt_T [1] ), .QN(_103_ ) );
DFF_X1 \g_mem.delayCnt_prng.state_2_$_SDFF_PP0__Q ( .D(_042_ ), .CK(clock ), .Q(\g_mem._delayCnt_T [2] ), .QN(_102_ ) );
DFF_X1 \g_mem.mem_data_Reg_$_SDFFE_PP0P__Q ( .D(_004_ ), .CK(_096_ ), .Q(\c_arbiter.io_axi_r_data [2] ), .QN(_139_ ) );
DFF_X1 \g_mem.mem_data_Reg_$_SDFFE_PP0P__Q_1 ( .D(_043_ ), .CK(_096_ ), .Q(\c_arbiter.io_axi_r_data [1] ), .QN(_101_ ) );
DFF_X1 \g_mem.mem_data_Reg_$_SDFFE_PP0P__Q_2 ( .D(_044_ ), .CK(_096_ ), .Q(\c_arbiter.io_axi_r_data [0] ), .QN(_100_ ) );
DFF_X1 \g_mem.validReg_$_SDFF_PP0__Q ( .D(_045_ ), .CK(clock ), .Q(\g_mem.validReg ), .QN(_099_ ) );

endmodule
