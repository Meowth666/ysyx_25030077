//Generate the verilog at 2025-05-25T16:24:40 by iSTA.
module MyOperators (
clk,
io_carry,
io_overflow,
reset,
io_in_a,
io_in_b,
io_out,
io_sw
);

input clk ;
output io_carry ;
output io_overflow ;
input reset ;
input [31:0] io_in_a ;
input [31:0] io_in_b ;
output [31:0] io_out ;
input [3:0] io_sw ;

wire _0000_ ;
wire _0001_ ;
wire _0002_ ;
wire _0003_ ;
wire _0004_ ;
wire _0005_ ;
wire _0006_ ;
wire _0007_ ;
wire _0008_ ;
wire _0009_ ;
wire _0010_ ;
wire _0011_ ;
wire _0012_ ;
wire _0013_ ;
wire _0014_ ;
wire _0015_ ;
wire _0016_ ;
wire _0017_ ;
wire _0018_ ;
wire _0019_ ;
wire _0020_ ;
wire _0021_ ;
wire _0022_ ;
wire _0023_ ;
wire _0024_ ;
wire _0025_ ;
wire _0026_ ;
wire _0027_ ;
wire _0028_ ;
wire _0029_ ;
wire _0030_ ;
wire _0031_ ;
wire _0032_ ;
wire _0033_ ;
wire _0034_ ;
wire _0035_ ;
wire _0036_ ;
wire _0037_ ;
wire _0038_ ;
wire _0039_ ;
wire _0040_ ;
wire _0041_ ;
wire _0042_ ;
wire _0043_ ;
wire _0044_ ;
wire _0045_ ;
wire _0046_ ;
wire _0047_ ;
wire _0048_ ;
wire _0049_ ;
wire _0050_ ;
wire _0051_ ;
wire _0052_ ;
wire _0053_ ;
wire _0054_ ;
wire _0055_ ;
wire _0056_ ;
wire _0057_ ;
wire _0058_ ;
wire _0059_ ;
wire _0060_ ;
wire _0061_ ;
wire _0062_ ;
wire _0063_ ;
wire _0064_ ;
wire _0065_ ;
wire _0066_ ;
wire _0067_ ;
wire _0068_ ;
wire _0069_ ;
wire _0070_ ;
wire _0071_ ;
wire _0072_ ;
wire _0073_ ;
wire _0074_ ;
wire _0075_ ;
wire _0076_ ;
wire _0077_ ;
wire _0078_ ;
wire _0079_ ;
wire _0080_ ;
wire _0081_ ;
wire _0082_ ;
wire _0083_ ;
wire _0084_ ;
wire _0085_ ;
wire _0086_ ;
wire _0087_ ;
wire _0088_ ;
wire _0089_ ;
wire _0090_ ;
wire _0091_ ;
wire _0092_ ;
wire _0093_ ;
wire _0094_ ;
wire _0095_ ;
wire _0096_ ;
wire _0097_ ;
wire _0098_ ;
wire _0099_ ;
wire _0100_ ;
wire _0101_ ;
wire _0102_ ;
wire _0103_ ;
wire _0104_ ;
wire _0105_ ;
wire _0106_ ;
wire _0107_ ;
wire _0108_ ;
wire _0109_ ;
wire _0110_ ;
wire _0111_ ;
wire _0112_ ;
wire _0113_ ;
wire _0114_ ;
wire _0115_ ;
wire _0116_ ;
wire _0117_ ;
wire _0118_ ;
wire _0119_ ;
wire _0120_ ;
wire _0121_ ;
wire _0122_ ;
wire _0123_ ;
wire _0124_ ;
wire _0125_ ;
wire _0126_ ;
wire _0127_ ;
wire _0128_ ;
wire _0129_ ;
wire _0130_ ;
wire _0131_ ;
wire _0132_ ;
wire _0133_ ;
wire _0134_ ;
wire _0135_ ;
wire _0136_ ;
wire _0137_ ;
wire _0138_ ;
wire _0139_ ;
wire _0140_ ;
wire _0141_ ;
wire _0142_ ;
wire _0143_ ;
wire _0144_ ;
wire _0145_ ;
wire _0146_ ;
wire _0147_ ;
wire _0148_ ;
wire _0149_ ;
wire _0150_ ;
wire _0151_ ;
wire _0152_ ;
wire _0153_ ;
wire _0154_ ;
wire _0155_ ;
wire _0156_ ;
wire _0157_ ;
wire _0158_ ;
wire _0159_ ;
wire _0160_ ;
wire _0161_ ;
wire _0162_ ;
wire _0163_ ;
wire _0164_ ;
wire _0165_ ;
wire _0166_ ;
wire _0167_ ;
wire _0168_ ;
wire _0169_ ;
wire _0170_ ;
wire _0171_ ;
wire _0172_ ;
wire _0173_ ;
wire _0174_ ;
wire _0175_ ;
wire _0176_ ;
wire _0177_ ;
wire _0178_ ;
wire _0179_ ;
wire _0180_ ;
wire _0181_ ;
wire _0182_ ;
wire _0183_ ;
wire _0184_ ;
wire _0185_ ;
wire _0186_ ;
wire _0187_ ;
wire _0188_ ;
wire _0189_ ;
wire _0190_ ;
wire _0191_ ;
wire _0192_ ;
wire _0193_ ;
wire _0194_ ;
wire _0195_ ;
wire _0196_ ;
wire _0197_ ;
wire _0198_ ;
wire _0199_ ;
wire _0200_ ;
wire _0201_ ;
wire _0202_ ;
wire _0203_ ;
wire _0204_ ;
wire _0205_ ;
wire _0206_ ;
wire _0207_ ;
wire _0208_ ;
wire _0209_ ;
wire _0210_ ;
wire _0211_ ;
wire _0212_ ;
wire _0213_ ;
wire _0214_ ;
wire _0215_ ;
wire _0216_ ;
wire _0217_ ;
wire _0218_ ;
wire _0219_ ;
wire _0220_ ;
wire _0221_ ;
wire _0222_ ;
wire _0223_ ;
wire _0224_ ;
wire _0225_ ;
wire _0226_ ;
wire _0227_ ;
wire _0228_ ;
wire _0229_ ;
wire _0230_ ;
wire _0231_ ;
wire _0232_ ;
wire _0233_ ;
wire _0234_ ;
wire _0235_ ;
wire _0236_ ;
wire _0237_ ;
wire _0238_ ;
wire _0239_ ;
wire _0240_ ;
wire _0241_ ;
wire _0242_ ;
wire _0243_ ;
wire _0244_ ;
wire _0245_ ;
wire _0246_ ;
wire _0247_ ;
wire _0248_ ;
wire _0249_ ;
wire _0250_ ;
wire _0251_ ;
wire _0252_ ;
wire _0253_ ;
wire _0254_ ;
wire _0255_ ;
wire _0256_ ;
wire _0257_ ;
wire _0258_ ;
wire _0259_ ;
wire _0260_ ;
wire _0261_ ;
wire _0262_ ;
wire _0263_ ;
wire _0264_ ;
wire _0265_ ;
wire _0266_ ;
wire _0267_ ;
wire _0268_ ;
wire _0269_ ;
wire _0270_ ;
wire _0271_ ;
wire _0272_ ;
wire _0273_ ;
wire _0274_ ;
wire _0275_ ;
wire _0276_ ;
wire _0277_ ;
wire _0278_ ;
wire _0279_ ;
wire _0280_ ;
wire _0281_ ;
wire _0282_ ;
wire _0283_ ;
wire _0284_ ;
wire _0285_ ;
wire _0286_ ;
wire _0287_ ;
wire _0288_ ;
wire _0289_ ;
wire _0290_ ;
wire _0291_ ;
wire _0292_ ;
wire _0293_ ;
wire _0294_ ;
wire _0295_ ;
wire _0296_ ;
wire _0297_ ;
wire _0298_ ;
wire _0299_ ;
wire _0300_ ;
wire _0301_ ;
wire _0302_ ;
wire _0303_ ;
wire _0304_ ;
wire _0305_ ;
wire _0306_ ;
wire _0307_ ;
wire _0308_ ;
wire _0309_ ;
wire _0310_ ;
wire _0311_ ;
wire _0312_ ;
wire _0313_ ;
wire _0314_ ;
wire _0315_ ;
wire _0316_ ;
wire _0317_ ;
wire _0318_ ;
wire _0319_ ;
wire _0320_ ;
wire _0321_ ;
wire _0322_ ;
wire _0323_ ;
wire _0324_ ;
wire _0325_ ;
wire _0326_ ;
wire _0327_ ;
wire _0328_ ;
wire _0329_ ;
wire _0330_ ;
wire _0331_ ;
wire _0332_ ;
wire _0333_ ;
wire _0334_ ;
wire _0335_ ;
wire _0336_ ;
wire _0337_ ;
wire _0338_ ;
wire _0339_ ;
wire _0340_ ;
wire _0341_ ;
wire _0342_ ;
wire _0343_ ;
wire _0344_ ;
wire _0345_ ;
wire _0346_ ;
wire _0347_ ;
wire _0348_ ;
wire _0349_ ;
wire _0350_ ;
wire _0351_ ;
wire _0352_ ;
wire _0353_ ;
wire _0354_ ;
wire _0355_ ;
wire _0356_ ;
wire _0357_ ;
wire _0358_ ;
wire _0359_ ;
wire _0360_ ;
wire _0361_ ;
wire _0362_ ;
wire _0363_ ;
wire _0364_ ;
wire _0365_ ;
wire _0366_ ;
wire _0367_ ;
wire _0368_ ;
wire _0369_ ;
wire _0370_ ;
wire _0371_ ;
wire _0372_ ;
wire _0373_ ;
wire _0374_ ;
wire _0375_ ;
wire _0376_ ;
wire _0377_ ;
wire _0378_ ;
wire _0379_ ;
wire _0380_ ;
wire _0381_ ;
wire _0382_ ;
wire _0383_ ;
wire _0384_ ;
wire _0385_ ;
wire _0386_ ;
wire _0387_ ;
wire _0388_ ;
wire _0389_ ;
wire _0390_ ;
wire _0391_ ;
wire _0392_ ;
wire _0393_ ;
wire _0394_ ;
wire _0395_ ;
wire _0396_ ;
wire _0397_ ;
wire _0398_ ;
wire _0399_ ;
wire _0400_ ;
wire _0401_ ;
wire _0402_ ;
wire _0403_ ;
wire _0404_ ;
wire _0405_ ;
wire _0406_ ;
wire _0407_ ;
wire _0408_ ;
wire _0409_ ;
wire _0410_ ;
wire _0411_ ;
wire _0412_ ;
wire _0413_ ;
wire _0414_ ;
wire _0415_ ;
wire _0416_ ;
wire _0417_ ;
wire _0418_ ;
wire _0419_ ;
wire _0420_ ;
wire _0421_ ;
wire _0422_ ;
wire _0423_ ;
wire _0424_ ;
wire _0425_ ;
wire _0426_ ;
wire _0427_ ;
wire _0428_ ;
wire _0429_ ;
wire _0430_ ;
wire _0431_ ;
wire _0432_ ;
wire _0433_ ;
wire _0434_ ;
wire _0435_ ;
wire _0436_ ;
wire _0437_ ;
wire _0438_ ;
wire _0439_ ;
wire _0440_ ;
wire _0441_ ;
wire _0442_ ;
wire _0443_ ;
wire _0444_ ;
wire _0445_ ;
wire _0446_ ;
wire _0447_ ;
wire _0448_ ;
wire _0449_ ;
wire _0450_ ;
wire _0451_ ;
wire _0452_ ;
wire _0453_ ;
wire _0454_ ;
wire _0455_ ;
wire _0456_ ;
wire _0457_ ;
wire _0458_ ;
wire _0459_ ;
wire _0460_ ;
wire _0461_ ;
wire _0462_ ;
wire _0463_ ;
wire _0464_ ;
wire _0465_ ;
wire _0466_ ;
wire _0467_ ;
wire _0468_ ;
wire _0469_ ;
wire _0470_ ;
wire _0471_ ;
wire _0472_ ;
wire _0473_ ;
wire _0474_ ;
wire _0475_ ;
wire _0476_ ;
wire _0477_ ;
wire _0478_ ;
wire _0479_ ;
wire _0480_ ;
wire _0481_ ;
wire _0482_ ;
wire _0483_ ;
wire _0484_ ;
wire _0485_ ;
wire _0486_ ;
wire _0487_ ;
wire _0488_ ;
wire _0489_ ;
wire _0490_ ;
wire _0491_ ;
wire _0492_ ;
wire _0493_ ;
wire _0494_ ;
wire _0495_ ;
wire _0496_ ;
wire _0497_ ;
wire _0498_ ;
wire _0499_ ;
wire _0500_ ;
wire _0501_ ;
wire _0502_ ;
wire _0503_ ;
wire _0504_ ;
wire _0505_ ;
wire _0506_ ;
wire _0507_ ;
wire _0508_ ;
wire _0509_ ;
wire _0510_ ;
wire _0511_ ;
wire _0512_ ;
wire _0513_ ;
wire _0514_ ;
wire _0515_ ;
wire _0516_ ;
wire _0517_ ;
wire _0518_ ;
wire _0519_ ;
wire _0520_ ;
wire _0521_ ;
wire _0522_ ;
wire _0523_ ;
wire _0524_ ;
wire _0525_ ;
wire _0526_ ;
wire _0527_ ;
wire _0528_ ;
wire _0529_ ;
wire _0530_ ;
wire _0531_ ;
wire _0532_ ;
wire _0533_ ;
wire _0534_ ;
wire _0535_ ;
wire _0536_ ;
wire _0537_ ;
wire _0538_ ;
wire _0539_ ;
wire _0540_ ;
wire _0541_ ;
wire _0542_ ;
wire _0543_ ;
wire _0544_ ;
wire _0545_ ;
wire _0546_ ;
wire _0547_ ;
wire _0548_ ;
wire _0549_ ;
wire _0550_ ;
wire _0551_ ;
wire _0552_ ;
wire _0553_ ;
wire _0554_ ;
wire _0555_ ;
wire _0556_ ;
wire _0557_ ;
wire _0558_ ;
wire _0559_ ;
wire _0560_ ;
wire _0561_ ;
wire _0562_ ;
wire _0563_ ;
wire _0564_ ;
wire _0565_ ;
wire _0566_ ;
wire _0567_ ;
wire _0568_ ;
wire _0569_ ;
wire _0570_ ;
wire _0571_ ;
wire _0572_ ;
wire _0573_ ;
wire _0574_ ;
wire _0575_ ;
wire _0576_ ;
wire _0577_ ;
wire _0578_ ;
wire _0579_ ;
wire _0580_ ;
wire _0581_ ;
wire _0582_ ;
wire _0583_ ;
wire _0584_ ;
wire _0585_ ;
wire _0586_ ;
wire _0587_ ;
wire _0588_ ;
wire _0589_ ;
wire _0590_ ;
wire _0591_ ;
wire _0592_ ;
wire _0593_ ;
wire _0594_ ;
wire _0595_ ;
wire _0596_ ;
wire _0597_ ;
wire _0598_ ;
wire _0599_ ;
wire _0600_ ;
wire _0601_ ;
wire _0602_ ;
wire _0603_ ;
wire _0604_ ;
wire _0605_ ;
wire _0606_ ;
wire _0607_ ;
wire _0608_ ;
wire _0609_ ;
wire _0610_ ;
wire _0611_ ;
wire _0612_ ;
wire _0613_ ;
wire _0614_ ;
wire _0615_ ;
wire _0616_ ;
wire _0617_ ;
wire _0618_ ;
wire _0619_ ;
wire _0620_ ;
wire _0621_ ;
wire _0622_ ;
wire _0623_ ;
wire _0624_ ;
wire _0625_ ;
wire _0626_ ;
wire _0627_ ;
wire _0628_ ;
wire _0629_ ;
wire _0630_ ;
wire _0631_ ;
wire _0632_ ;
wire _0633_ ;
wire _0634_ ;
wire _0635_ ;
wire _0636_ ;
wire _0637_ ;
wire _0638_ ;
wire _0639_ ;
wire _0640_ ;
wire _0641_ ;
wire _0642_ ;
wire _0643_ ;
wire _0644_ ;
wire _0645_ ;
wire _0646_ ;
wire _0647_ ;
wire _0648_ ;
wire _0649_ ;
wire _0650_ ;
wire _0651_ ;
wire _0652_ ;
wire _0653_ ;
wire _0654_ ;
wire _0655_ ;
wire _0656_ ;
wire _0657_ ;
wire _0658_ ;
wire _0659_ ;
wire _0660_ ;
wire _0661_ ;
wire _0662_ ;
wire _0663_ ;
wire _0664_ ;
wire _0665_ ;
wire _0666_ ;
wire _0667_ ;
wire _0668_ ;
wire _0669_ ;
wire _0670_ ;
wire _0671_ ;
wire _0672_ ;
wire _0673_ ;
wire _0674_ ;
wire _0675_ ;
wire _0676_ ;
wire _0677_ ;
wire _0678_ ;
wire _0679_ ;
wire _0680_ ;
wire _0681_ ;
wire _0682_ ;
wire _0683_ ;
wire _0684_ ;
wire _0685_ ;
wire _0686_ ;
wire _0687_ ;
wire _0688_ ;
wire _0689_ ;
wire _0690_ ;
wire _0691_ ;
wire _0692_ ;
wire _0693_ ;
wire _0694_ ;
wire _0695_ ;
wire _0696_ ;
wire _0697_ ;
wire _0698_ ;
wire _0699_ ;
wire _0700_ ;
wire _0701_ ;
wire _0702_ ;
wire _0703_ ;
wire _0704_ ;
wire _0705_ ;
wire _0706_ ;
wire _0707_ ;
wire _0708_ ;
wire _0709_ ;
wire _0710_ ;
wire _0711_ ;
wire _0712_ ;
wire _0713_ ;
wire _0714_ ;
wire _0715_ ;
wire _0716_ ;
wire _0717_ ;
wire _0718_ ;
wire _0719_ ;
wire _0720_ ;
wire _0721_ ;
wire _0722_ ;
wire _0723_ ;
wire _0724_ ;
wire _0725_ ;
wire _0726_ ;
wire _0727_ ;
wire _0728_ ;
wire _0729_ ;
wire _0730_ ;
wire _0731_ ;
wire _0732_ ;
wire _0733_ ;
wire _0734_ ;
wire _0735_ ;
wire _0736_ ;
wire _0737_ ;
wire _0738_ ;
wire _0739_ ;
wire _0740_ ;
wire _0741_ ;
wire _0742_ ;
wire _0743_ ;
wire _0744_ ;
wire _0745_ ;
wire _0746_ ;
wire _0747_ ;
wire _0748_ ;
wire _0749_ ;
wire _0750_ ;
wire _0751_ ;
wire _0752_ ;
wire _0753_ ;
wire _0754_ ;
wire _0755_ ;
wire _0756_ ;
wire _0757_ ;
wire _0758_ ;
wire _0759_ ;
wire _0760_ ;
wire _0761_ ;
wire _0762_ ;
wire _0763_ ;
wire _0764_ ;
wire _0765_ ;
wire _0766_ ;
wire _0767_ ;
wire _0768_ ;
wire _0769_ ;
wire _0770_ ;
wire _0771_ ;
wire _0772_ ;
wire _0773_ ;
wire _0774_ ;
wire _0775_ ;
wire _0776_ ;
wire _0777_ ;
wire _0778_ ;
wire _0779_ ;
wire _0780_ ;
wire _0781_ ;
wire _0782_ ;
wire _0783_ ;
wire _0784_ ;
wire _0785_ ;
wire _0786_ ;
wire _0787_ ;
wire _0788_ ;
wire _0789_ ;
wire _0790_ ;
wire _0791_ ;
wire _0792_ ;
wire _0793_ ;
wire _0794_ ;
wire _0795_ ;
wire _0796_ ;
wire _0797_ ;
wire _0798_ ;
wire _0799_ ;
wire _0800_ ;
wire _0801_ ;
wire _0802_ ;
wire _0803_ ;
wire _0804_ ;
wire _0805_ ;
wire _0806_ ;
wire _0807_ ;
wire _0808_ ;
wire _0809_ ;
wire _0810_ ;
wire _0811_ ;
wire _0812_ ;
wire _0813_ ;
wire _0814_ ;
wire _0815_ ;
wire _0816_ ;
wire _0817_ ;
wire _0818_ ;
wire _0819_ ;
wire _0820_ ;
wire _0821_ ;
wire _0822_ ;
wire _0823_ ;
wire _0824_ ;
wire _0825_ ;
wire _0826_ ;
wire _0827_ ;
wire _0828_ ;
wire _0829_ ;
wire _0830_ ;
wire _0831_ ;
wire _0832_ ;
wire _0833_ ;
wire _0834_ ;
wire _0835_ ;
wire _0836_ ;
wire _0837_ ;
wire _0838_ ;
wire _0839_ ;
wire _0840_ ;
wire _0841_ ;
wire _0842_ ;
wire _0843_ ;
wire _0844_ ;
wire _0845_ ;
wire _0846_ ;
wire _0847_ ;
wire _0848_ ;
wire _0849_ ;
wire _0850_ ;
wire _0851_ ;
wire _0852_ ;
wire _0853_ ;
wire _0854_ ;
wire _0855_ ;
wire _0856_ ;
wire _0857_ ;
wire _0858_ ;
wire _0859_ ;
wire _0860_ ;
wire _0861_ ;
wire _0862_ ;
wire _0863_ ;
wire _0864_ ;
wire _0865_ ;
wire _0866_ ;
wire _0867_ ;
wire _0868_ ;
wire _0869_ ;
wire _0870_ ;
wire _0871_ ;
wire _0872_ ;
wire _0873_ ;
wire _0874_ ;
wire _0875_ ;
wire _0876_ ;
wire _0877_ ;
wire _0878_ ;
wire _0879_ ;
wire _0880_ ;
wire _0881_ ;
wire _0882_ ;
wire _0883_ ;
wire _0884_ ;
wire _0885_ ;
wire _0886_ ;
wire _0887_ ;
wire _0888_ ;
wire _0889_ ;
wire _0890_ ;
wire _0891_ ;
wire _0892_ ;
wire _0893_ ;
wire _0894_ ;
wire _0895_ ;
wire _0896_ ;
wire _0897_ ;
wire _0898_ ;
wire _0899_ ;
wire _0900_ ;
wire _0901_ ;
wire _0902_ ;
wire _0903_ ;
wire _0904_ ;
wire _0905_ ;
wire _0906_ ;
wire _0907_ ;
wire _0908_ ;
wire _0909_ ;
wire _0910_ ;
wire _0911_ ;
wire _0912_ ;
wire _0913_ ;
wire _0914_ ;
wire _0915_ ;
wire _0916_ ;
wire _0917_ ;
wire _0918_ ;
wire _0919_ ;
wire _0920_ ;
wire _0921_ ;
wire _0922_ ;
wire _0923_ ;
wire _0924_ ;
wire _0925_ ;
wire _0926_ ;
wire _0927_ ;
wire _0928_ ;
wire _0929_ ;
wire _0930_ ;
wire _0931_ ;
wire _0932_ ;
wire _0933_ ;
wire _0934_ ;
wire _0935_ ;
wire _0936_ ;
wire _0937_ ;
wire _0938_ ;
wire _0939_ ;
wire _0940_ ;
wire _0941_ ;
wire _0942_ ;
wire _0943_ ;
wire _0944_ ;
wire _0945_ ;
wire _0946_ ;
wire _0947_ ;
wire _0948_ ;
wire _0949_ ;
wire _0950_ ;
wire _0951_ ;
wire _0952_ ;
wire _0953_ ;
wire _0954_ ;
wire _0955_ ;
wire _0956_ ;
wire _0957_ ;
wire _0958_ ;
wire _0959_ ;
wire _0960_ ;
wire _0961_ ;
wire _0962_ ;
wire _0963_ ;
wire _0964_ ;
wire _0965_ ;
wire _0966_ ;
wire _0967_ ;
wire _0968_ ;
wire _0969_ ;
wire _0970_ ;
wire _0971_ ;
wire _0972_ ;
wire _0973_ ;
wire _0974_ ;
wire _0975_ ;
wire _0976_ ;
wire _0977_ ;
wire _0978_ ;
wire _0979_ ;
wire _0980_ ;
wire _0981_ ;
wire _0982_ ;
wire _0983_ ;
wire _0984_ ;
wire _0985_ ;
wire _0986_ ;
wire _0987_ ;
wire _0988_ ;
wire _0989_ ;
wire _0990_ ;
wire _0991_ ;
wire _0992_ ;
wire _0993_ ;
wire _0994_ ;
wire _0995_ ;
wire _0996_ ;
wire _0997_ ;
wire _0998_ ;
wire _0999_ ;
wire _1000_ ;
wire _1001_ ;
wire _1002_ ;
wire _1003_ ;
wire _1004_ ;
wire _1005_ ;
wire _1006_ ;
wire _1007_ ;
wire _1008_ ;
wire _1009_ ;
wire _1010_ ;
wire _1011_ ;
wire _1012_ ;
wire _1013_ ;
wire _1014_ ;
wire _1015_ ;
wire _1016_ ;
wire _1017_ ;
wire _1018_ ;
wire _1019_ ;
wire _1020_ ;
wire _1021_ ;
wire _1022_ ;
wire _1023_ ;
wire _1024_ ;
wire _1025_ ;
wire _1026_ ;
wire _1027_ ;
wire _1028_ ;
wire _1029_ ;
wire _1030_ ;
wire _1031_ ;
wire _1032_ ;
wire _1033_ ;
wire _1034_ ;
wire _1035_ ;
wire _1036_ ;
wire _1037_ ;
wire _1038_ ;
wire _1039_ ;
wire _1040_ ;
wire _1041_ ;
wire _1042_ ;
wire _1043_ ;
wire _1044_ ;
wire _1045_ ;
wire _1046_ ;
wire _1047_ ;
wire _1048_ ;
wire _1049_ ;
wire _1050_ ;
wire _1051_ ;
wire _1052_ ;
wire _1053_ ;
wire _1054_ ;
wire _1055_ ;
wire _1056_ ;
wire _1057_ ;
wire _1058_ ;
wire _1059_ ;
wire _1060_ ;
wire _1061_ ;
wire _1062_ ;
wire _1063_ ;
wire _1064_ ;
wire _1065_ ;
wire _1066_ ;
wire _1067_ ;
wire _1068_ ;
wire _1069_ ;
wire _1070_ ;
wire _1071_ ;
wire _1072_ ;
wire _1073_ ;
wire _1074_ ;
wire _1075_ ;
wire _1076_ ;
wire _1077_ ;
wire _1078_ ;
wire _1079_ ;
wire _1080_ ;
wire _1081_ ;
wire _1082_ ;
wire _1083_ ;
wire _1084_ ;
wire _1085_ ;
wire _1086_ ;
wire _1087_ ;
wire _1088_ ;
wire _1089_ ;
wire _1090_ ;
wire _1091_ ;
wire _1092_ ;
wire _1093_ ;
wire _1094_ ;
wire _1095_ ;
wire _1096_ ;
wire _1097_ ;
wire _1098_ ;
wire _1099_ ;
wire _1100_ ;
wire _1101_ ;
wire _1102_ ;
wire _1103_ ;
wire _1104_ ;
wire _1105_ ;
wire _1106_ ;
wire _1107_ ;
wire _1108_ ;
wire _1109_ ;
wire _1110_ ;
wire _1111_ ;
wire _1112_ ;
wire _1113_ ;
wire _1114_ ;
wire _1115_ ;
wire _1116_ ;
wire _1117_ ;
wire _1118_ ;
wire _1119_ ;
wire _1120_ ;
wire _1121_ ;
wire _1122_ ;
wire _1123_ ;
wire _1124_ ;
wire _1125_ ;
wire _1126_ ;
wire _1127_ ;
wire _1128_ ;
wire _1129_ ;
wire _1130_ ;
wire _1131_ ;
wire _1132_ ;
wire _1133_ ;
wire _1134_ ;
wire _1135_ ;
wire _1136_ ;
wire _1137_ ;
wire _1138_ ;
wire _1139_ ;
wire _1140_ ;
wire _1141_ ;
wire _1142_ ;
wire _1143_ ;
wire _1144_ ;
wire _1145_ ;
wire _1146_ ;
wire _1147_ ;
wire _1148_ ;
wire _1149_ ;
wire _1150_ ;
wire _1151_ ;
wire _1152_ ;
wire _1153_ ;
wire _1154_ ;
wire _1155_ ;
wire _1156_ ;
wire _1157_ ;
wire _1158_ ;
wire _1159_ ;
wire _1160_ ;
wire _1161_ ;
wire _1162_ ;
wire _1163_ ;
wire _1164_ ;
wire _1165_ ;
wire _1166_ ;
wire _1167_ ;
wire _1168_ ;
wire _1169_ ;
wire _1170_ ;
wire _1171_ ;
wire _1172_ ;
wire _1173_ ;
wire _1174_ ;
wire _1175_ ;
wire _1176_ ;
wire _1177_ ;
wire _1178_ ;
wire _1179_ ;
wire _1180_ ;
wire _1181_ ;
wire _1182_ ;
wire _1183_ ;
wire _1184_ ;
wire _1185_ ;
wire _1186_ ;
wire _1187_ ;
wire _1188_ ;
wire _1189_ ;
wire _1190_ ;
wire _1191_ ;
wire _1192_ ;
wire _1193_ ;
wire _1194_ ;
wire _1195_ ;
wire _1196_ ;
wire _1197_ ;
wire _1198_ ;
wire _1199_ ;
wire _1200_ ;
wire _1201_ ;
wire _1202_ ;
wire _1203_ ;
wire _1204_ ;
wire _1205_ ;
wire _1206_ ;
wire _1207_ ;
wire _1208_ ;
wire _1209_ ;
wire _1210_ ;
wire _1211_ ;
wire _1212_ ;
wire _1213_ ;
wire _1214_ ;
wire _1215_ ;
wire _1216_ ;
wire _1217_ ;
wire _1218_ ;
wire _1219_ ;
wire _1220_ ;
wire _1221_ ;
wire _1222_ ;
wire _1223_ ;
wire _1224_ ;
wire _1225_ ;
wire _1226_ ;
wire _1227_ ;
wire _1228_ ;
wire _1229_ ;
wire _1230_ ;
wire _1231_ ;
wire _1232_ ;
wire _1233_ ;
wire _1234_ ;
wire _1235_ ;
wire _1236_ ;
wire _1237_ ;
wire _1238_ ;
wire _1239_ ;
wire _1240_ ;
wire _1241_ ;
wire _1242_ ;
wire _1243_ ;
wire _1244_ ;
wire _1245_ ;
wire _1246_ ;
wire _1247_ ;
wire _1248_ ;
wire _1249_ ;
wire _1250_ ;
wire _1251_ ;
wire _1252_ ;
wire _1253_ ;
wire _1254_ ;
wire _1255_ ;
wire _1256_ ;
wire _1257_ ;
wire _1258_ ;
wire _1259_ ;
wire _1260_ ;
wire _1261_ ;
wire _1262_ ;
wire _1263_ ;
wire _1264_ ;
wire _1265_ ;
wire _1266_ ;
wire _1267_ ;
wire _1268_ ;
wire _1269_ ;
wire _1270_ ;
wire _1271_ ;
wire _1272_ ;
wire _1273_ ;
wire _1274_ ;
wire _1275_ ;
wire _1276_ ;
wire _1277_ ;
wire _1278_ ;
wire _1279_ ;
wire _1280_ ;
wire _1281_ ;
wire _1282_ ;
wire _1283_ ;
wire _1284_ ;
wire _1285_ ;
wire _1286_ ;
wire _1287_ ;
wire _1288_ ;
wire _1289_ ;
wire _1290_ ;
wire _1291_ ;
wire _1292_ ;
wire _1293_ ;
wire _1294_ ;
wire _1295_ ;
wire _1296_ ;
wire _1297_ ;
wire _1298_ ;
wire _1299_ ;
wire _1300_ ;
wire _1301_ ;
wire _1302_ ;
wire _1303_ ;
wire _1304_ ;
wire _1305_ ;
wire _1306_ ;
wire _1307_ ;
wire _1308_ ;
wire _1309_ ;
wire _1310_ ;
wire _1311_ ;
wire _1312_ ;
wire _1313_ ;
wire _1314_ ;
wire _1315_ ;
wire _1316_ ;
wire _1317_ ;
wire _1318_ ;
wire _1319_ ;
wire _1320_ ;
wire _1321_ ;
wire _1322_ ;
wire _1323_ ;
wire _1324_ ;
wire _1325_ ;
wire _1326_ ;
wire _1327_ ;
wire _1328_ ;
wire _1329_ ;
wire _1330_ ;
wire _1331_ ;
wire _1332_ ;
wire _1333_ ;
wire _1334_ ;
wire _1335_ ;
wire _1336_ ;
wire _1337_ ;
wire _1338_ ;
wire _1339_ ;
wire _1340_ ;
wire _1341_ ;
wire _1342_ ;
wire _1343_ ;
wire _1344_ ;
wire _1345_ ;
wire _1346_ ;
wire _1347_ ;
wire _1348_ ;
wire _1349_ ;
wire _1350_ ;
wire _1351_ ;
wire _1352_ ;
wire _1353_ ;
wire _1354_ ;
wire _1355_ ;
wire _1356_ ;
wire _1357_ ;
wire _1358_ ;
wire _1359_ ;
wire _1360_ ;
wire _1361_ ;
wire _1362_ ;
wire _1363_ ;
wire _1364_ ;
wire _1365_ ;
wire _1366_ ;
wire _1367_ ;
wire _1368_ ;
wire _1369_ ;
wire _1370_ ;
wire _1371_ ;
wire _1372_ ;
wire _1373_ ;
wire _1374_ ;
wire _1375_ ;
wire _1376_ ;
wire _1377_ ;
wire _1378_ ;
wire _1379_ ;
wire _1380_ ;
wire _1381_ ;
wire _1382_ ;
wire _1383_ ;
wire _1384_ ;
wire _1385_ ;
wire _1386_ ;
wire _1387_ ;
wire _1388_ ;
wire _1389_ ;
wire _1390_ ;
wire _1391_ ;
wire _1392_ ;
wire _1393_ ;
wire _1394_ ;
wire _1395_ ;
wire _1396_ ;
wire _1397_ ;
wire _1398_ ;
wire _1399_ ;
wire _1400_ ;
wire _1401_ ;
wire _1402_ ;
wire _1403_ ;
wire _1404_ ;
wire _1405_ ;
wire _1406_ ;
wire _1407_ ;
wire _1408_ ;
wire _1409_ ;
wire _1410_ ;
wire _1411_ ;
wire _1412_ ;
wire _1413_ ;
wire _1414_ ;
wire _1415_ ;
wire _1416_ ;
wire _1417_ ;
wire _1418_ ;
wire _1419_ ;
wire _1420_ ;
wire _1421_ ;
wire _1422_ ;
wire _1423_ ;
wire _1424_ ;
wire _1425_ ;
wire _1426_ ;
wire _1427_ ;
wire _1428_ ;
wire _1429_ ;
wire _1430_ ;
wire _1431_ ;
wire _1432_ ;
wire _1433_ ;
wire _1434_ ;
wire _1435_ ;
wire _1436_ ;
wire _1437_ ;
wire _1438_ ;
wire _1439_ ;
wire _1440_ ;
wire _1441_ ;
wire _1442_ ;
wire _1443_ ;
wire _1444_ ;
wire _1445_ ;
wire _1446_ ;
wire _1447_ ;
wire _1448_ ;
wire _1449_ ;
wire _1450_ ;
wire _1451_ ;
wire _1452_ ;
wire _1453_ ;
wire _1454_ ;
wire _1455_ ;
wire _1456_ ;
wire _1457_ ;
wire _1458_ ;
wire _1459_ ;
wire _1460_ ;
wire _1461_ ;
wire _1462_ ;
wire _1463_ ;
wire _1464_ ;
wire _1465_ ;
wire _1466_ ;
wire _1467_ ;
wire _1468_ ;
wire _1469_ ;
wire _1470_ ;
wire _1471_ ;
wire _1472_ ;
wire _1473_ ;
wire _1474_ ;
wire _1475_ ;
wire _1476_ ;
wire _1477_ ;
wire _1478_ ;
wire _1479_ ;
wire _1480_ ;
wire _1481_ ;
wire _1482_ ;
wire _1483_ ;
wire _1484_ ;
wire _1485_ ;
wire _1486_ ;
wire _1487_ ;
wire _1488_ ;
wire _1489_ ;
wire _1490_ ;
wire _1491_ ;
wire _1492_ ;
wire _1493_ ;
wire _1494_ ;
wire _1495_ ;
wire _1496_ ;
wire _1497_ ;
wire _1498_ ;
wire _1499_ ;
wire _1500_ ;
wire _1501_ ;
wire _1502_ ;
wire _1503_ ;
wire _1504_ ;
wire _1505_ ;
wire _1506_ ;
wire _1507_ ;
wire _1508_ ;
wire _1509_ ;
wire _1510_ ;
wire _1511_ ;
wire _1512_ ;
wire _1513_ ;
wire _1514_ ;
wire _1515_ ;
wire _1516_ ;
wire _1517_ ;
wire _1518_ ;
wire _1519_ ;
wire _1520_ ;
wire _1521_ ;
wire _1522_ ;
wire _1523_ ;
wire _1524_ ;
wire _1525_ ;
wire _1526_ ;
wire _1527_ ;
wire _1528_ ;
wire _1529_ ;
wire _1530_ ;
wire _1531_ ;
wire _1532_ ;
wire _1533_ ;
wire _1534_ ;
wire _1535_ ;
wire _1536_ ;
wire _1537_ ;
wire _1538_ ;
wire _1539_ ;
wire _1540_ ;
wire _1541_ ;
wire _1542_ ;
wire _1543_ ;
wire _1544_ ;
wire _1545_ ;
wire _1546_ ;
wire _1547_ ;
wire _1548_ ;
wire _1549_ ;
wire _1550_ ;
wire _1551_ ;
wire _1552_ ;
wire _1553_ ;
wire _1554_ ;
wire _1555_ ;
wire _1556_ ;
wire _1557_ ;
wire _1558_ ;
wire _1559_ ;
wire _1560_ ;
wire _1561_ ;
wire _1562_ ;
wire _1563_ ;
wire _1564_ ;
wire _1565_ ;
wire _1566_ ;
wire _1567_ ;
wire _1568_ ;
wire _1569_ ;
wire _1570_ ;
wire _1571_ ;
wire _1572_ ;
wire _1573_ ;
wire _1574_ ;
wire _1575_ ;
wire _1576_ ;
wire _1577_ ;
wire _1578_ ;
wire _1579_ ;
wire _1580_ ;
wire _1581_ ;
wire _1582_ ;
wire _1583_ ;
wire _1584_ ;
wire _1585_ ;
wire _1586_ ;
wire _1587_ ;
wire _1588_ ;
wire _1589_ ;
wire _1590_ ;
wire _1591_ ;
wire _1592_ ;
wire _1593_ ;
wire _1594_ ;
wire _1595_ ;
wire _1596_ ;
wire _1597_ ;
wire _1598_ ;
wire _1599_ ;
wire _1600_ ;
wire _1601_ ;
wire _1602_ ;
wire _1603_ ;
wire _1604_ ;
wire _1605_ ;
wire _1606_ ;
wire _1607_ ;
wire _1608_ ;
wire _1609_ ;
wire _1610_ ;
wire _1611_ ;
wire _1612_ ;
wire _1613_ ;
wire _1614_ ;
wire _1615_ ;
wire _1616_ ;
wire _1617_ ;
wire _1618_ ;
wire _1619_ ;
wire _1620_ ;
wire _1621_ ;
wire _1622_ ;
wire _1623_ ;
wire _1624_ ;
wire _1625_ ;
wire _1626_ ;
wire _1627_ ;
wire _1628_ ;
wire _1629_ ;
wire _1630_ ;
wire _1631_ ;
wire _1632_ ;
wire _1633_ ;
wire _1634_ ;
wire _1635_ ;
wire _1636_ ;
wire _1637_ ;
wire _1638_ ;
wire _1639_ ;
wire _1640_ ;
wire _1641_ ;
wire _1642_ ;
wire _1643_ ;
wire _1644_ ;
wire _1645_ ;
wire _1646_ ;
wire _1647_ ;
wire _1648_ ;
wire _1649_ ;
wire _1650_ ;
wire _1651_ ;
wire _1652_ ;
wire _1653_ ;
wire _1654_ ;
wire _1655_ ;
wire _1656_ ;
wire _1657_ ;
wire _1658_ ;
wire _1659_ ;
wire _1660_ ;
wire _1661_ ;
wire _1662_ ;
wire _1663_ ;
wire _1664_ ;
wire _1665_ ;
wire _1666_ ;
wire _1667_ ;
wire _1668_ ;
wire _1669_ ;
wire _1670_ ;
wire _1671_ ;
wire _1672_ ;
wire _1673_ ;
wire _1674_ ;
wire _1675_ ;
wire _1676_ ;
wire _1677_ ;
wire _1678_ ;
wire _1679_ ;
wire _1680_ ;
wire _1681_ ;
wire _1682_ ;
wire _1683_ ;
wire _1684_ ;
wire _1685_ ;
wire _1686_ ;
wire _1687_ ;
wire _1688_ ;
wire _1689_ ;
wire _1690_ ;
wire _1691_ ;
wire _1692_ ;
wire _1693_ ;
wire _1694_ ;
wire _1695_ ;
wire _1696_ ;
wire _1697_ ;
wire _1698_ ;
wire _1699_ ;
wire _1700_ ;
wire _1701_ ;
wire _1702_ ;
wire _1703_ ;
wire _1704_ ;
wire _1705_ ;
wire _1706_ ;
wire _1707_ ;
wire _1708_ ;
wire _1709_ ;
wire _1710_ ;
wire _1711_ ;
wire _1712_ ;
wire _1713_ ;
wire _1714_ ;
wire _1715_ ;
wire _1716_ ;
wire _1717_ ;
wire _1718_ ;
wire _1719_ ;
wire _1720_ ;
wire _1721_ ;
wire _1722_ ;
wire _1723_ ;
wire _1724_ ;
wire _1725_ ;
wire _1726_ ;
wire _1727_ ;
wire _1728_ ;
wire _1729_ ;
wire _1730_ ;
wire _1731_ ;
wire _1732_ ;
wire _1733_ ;
wire _1734_ ;
wire _1735_ ;
wire _1736_ ;
wire _1737_ ;
wire _1738_ ;
wire _1739_ ;
wire _1740_ ;
wire _1741_ ;
wire _1742_ ;
wire _1743_ ;
wire _1744_ ;
wire _1745_ ;
wire _1746_ ;
wire _1747_ ;
wire _1748_ ;
wire _1749_ ;
wire _1750_ ;
wire _1751_ ;
wire _1752_ ;
wire _1753_ ;
wire _1754_ ;
wire _1755_ ;
wire _1756_ ;
wire _1757_ ;
wire _1758_ ;
wire _1759_ ;
wire _1760_ ;
wire _1761_ ;
wire _1762_ ;
wire _1763_ ;
wire _1764_ ;
wire _1765_ ;
wire _1766_ ;
wire _1767_ ;
wire _1768_ ;
wire _1769_ ;
wire _1770_ ;
wire _1771_ ;
wire _1772_ ;
wire _1773_ ;
wire _1774_ ;
wire _1775_ ;
wire _1776_ ;
wire _1777_ ;
wire _1778_ ;
wire _1779_ ;
wire _1780_ ;
wire _1781_ ;
wire _1782_ ;
wire _1783_ ;
wire _1784_ ;
wire _1785_ ;
wire _1786_ ;
wire _1787_ ;
wire _1788_ ;
wire _1789_ ;
wire _1790_ ;
wire _1791_ ;
wire _1792_ ;
wire _1793_ ;
wire _1794_ ;
wire _1795_ ;
wire _1796_ ;
wire _1797_ ;
wire _1798_ ;
wire _1799_ ;
wire _1800_ ;
wire _1801_ ;
wire _1802_ ;
wire _1803_ ;
wire _1804_ ;
wire _1805_ ;
wire _1806_ ;
wire _1807_ ;
wire _1808_ ;
wire _1809_ ;
wire _1810_ ;
wire clk ;
wire io_carry ;
wire io_overflow ;
wire reset ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire \io_in_a[0] ;
wire \io_in_a[1] ;
wire \io_in_a[2] ;
wire \io_in_a[3] ;
wire \io_in_a[4] ;
wire \io_in_a[5] ;
wire \io_in_a[6] ;
wire \io_in_a[7] ;
wire \io_in_a[8] ;
wire \io_in_a[9] ;
wire \io_in_a[10] ;
wire \io_in_a[11] ;
wire \io_in_a[12] ;
wire \io_in_a[13] ;
wire \io_in_a[14] ;
wire \io_in_a[15] ;
wire \io_in_a[16] ;
wire \io_in_a[17] ;
wire \io_in_a[18] ;
wire \io_in_a[19] ;
wire \io_in_a[20] ;
wire \io_in_a[21] ;
wire \io_in_a[22] ;
wire \io_in_a[23] ;
wire \io_in_a[24] ;
wire \io_in_a[25] ;
wire \io_in_a[26] ;
wire \io_in_a[27] ;
wire \io_in_a[28] ;
wire \io_in_a[29] ;
wire \io_in_a[30] ;
wire \io_in_a[31] ;
wire \io_in_b[0] ;
wire \io_in_b[1] ;
wire \io_in_b[2] ;
wire \io_in_b[3] ;
wire \io_in_b[4] ;
wire \io_in_b[5] ;
wire \io_in_b[6] ;
wire \io_in_b[7] ;
wire \io_in_b[8] ;
wire \io_in_b[9] ;
wire \io_in_b[10] ;
wire \io_in_b[11] ;
wire \io_in_b[12] ;
wire \io_in_b[13] ;
wire \io_in_b[14] ;
wire \io_in_b[15] ;
wire \io_in_b[16] ;
wire \io_in_b[17] ;
wire \io_in_b[18] ;
wire \io_in_b[19] ;
wire \io_in_b[20] ;
wire \io_in_b[21] ;
wire \io_in_b[22] ;
wire \io_in_b[23] ;
wire \io_in_b[24] ;
wire \io_in_b[25] ;
wire \io_in_b[26] ;
wire \io_in_b[27] ;
wire \io_in_b[28] ;
wire \io_in_b[29] ;
wire \io_in_b[30] ;
wire \io_in_b[31] ;
wire \io_out[0] ;
wire \io_out[1] ;
wire \io_out[2] ;
wire \io_out[3] ;
wire \io_out[4] ;
wire \io_out[5] ;
wire \io_out[6] ;
wire \io_out[7] ;
wire \io_out[8] ;
wire \io_out[9] ;
wire \io_out[10] ;
wire \io_out[11] ;
wire \io_out[12] ;
wire \io_out[13] ;
wire \io_out[14] ;
wire \io_out[15] ;
wire \io_out[16] ;
wire \io_out[17] ;
wire \io_out[18] ;
wire \io_out[19] ;
wire \io_out[20] ;
wire \io_out[21] ;
wire \io_out[22] ;
wire \io_out[23] ;
wire \io_out[24] ;
wire \io_out[25] ;
wire \io_out[26] ;
wire \io_out[27] ;
wire \io_out[28] ;
wire \io_out[29] ;
wire \io_out[30] ;
wire \io_out[31] ;
wire \io_sw[0] ;
wire \io_sw[1] ;
wire \io_sw[2] ;
wire \io_sw[3] ;

assign \io_in_a[0] = io_in_a[0] ;
assign \io_in_a[1] = io_in_a[1] ;
assign \io_in_a[2] = io_in_a[2] ;
assign \io_in_a[3] = io_in_a[3] ;
assign \io_in_a[4] = io_in_a[4] ;
assign \io_in_a[5] = io_in_a[5] ;
assign \io_in_a[6] = io_in_a[6] ;
assign \io_in_a[7] = io_in_a[7] ;
assign \io_in_a[8] = io_in_a[8] ;
assign \io_in_a[9] = io_in_a[9] ;
assign \io_in_a[10] = io_in_a[10] ;
assign \io_in_a[11] = io_in_a[11] ;
assign \io_in_a[12] = io_in_a[12] ;
assign \io_in_a[13] = io_in_a[13] ;
assign \io_in_a[14] = io_in_a[14] ;
assign \io_in_a[15] = io_in_a[15] ;
assign \io_in_a[16] = io_in_a[16] ;
assign \io_in_a[17] = io_in_a[17] ;
assign \io_in_a[18] = io_in_a[18] ;
assign \io_in_a[19] = io_in_a[19] ;
assign \io_in_a[20] = io_in_a[20] ;
assign \io_in_a[21] = io_in_a[21] ;
assign \io_in_a[22] = io_in_a[22] ;
assign \io_in_a[23] = io_in_a[23] ;
assign \io_in_a[24] = io_in_a[24] ;
assign \io_in_a[25] = io_in_a[25] ;
assign \io_in_a[26] = io_in_a[26] ;
assign \io_in_a[27] = io_in_a[27] ;
assign \io_in_a[28] = io_in_a[28] ;
assign \io_in_a[29] = io_in_a[29] ;
assign \io_in_a[30] = io_in_a[30] ;
assign \io_in_a[31] = io_in_a[31] ;
assign \io_in_b[0] = io_in_b[0] ;
assign \io_in_b[1] = io_in_b[1] ;
assign \io_in_b[2] = io_in_b[2] ;
assign \io_in_b[3] = io_in_b[3] ;
assign \io_in_b[4] = io_in_b[4] ;
assign \io_in_b[5] = io_in_b[5] ;
assign \io_in_b[6] = io_in_b[6] ;
assign \io_in_b[7] = io_in_b[7] ;
assign \io_in_b[8] = io_in_b[8] ;
assign \io_in_b[9] = io_in_b[9] ;
assign \io_in_b[10] = io_in_b[10] ;
assign \io_in_b[11] = io_in_b[11] ;
assign \io_in_b[12] = io_in_b[12] ;
assign \io_in_b[13] = io_in_b[13] ;
assign \io_in_b[14] = io_in_b[14] ;
assign \io_in_b[15] = io_in_b[15] ;
assign \io_in_b[16] = io_in_b[16] ;
assign \io_in_b[17] = io_in_b[17] ;
assign \io_in_b[18] = io_in_b[18] ;
assign \io_in_b[19] = io_in_b[19] ;
assign \io_in_b[20] = io_in_b[20] ;
assign \io_in_b[21] = io_in_b[21] ;
assign \io_in_b[22] = io_in_b[22] ;
assign \io_in_b[23] = io_in_b[23] ;
assign \io_in_b[24] = io_in_b[24] ;
assign \io_in_b[25] = io_in_b[25] ;
assign \io_in_b[26] = io_in_b[26] ;
assign \io_in_b[27] = io_in_b[27] ;
assign \io_in_b[28] = io_in_b[28] ;
assign \io_in_b[29] = io_in_b[29] ;
assign \io_in_b[30] = io_in_b[30] ;
assign \io_in_b[31] = io_in_b[31] ;
assign io_out[0] = \io_out[0] ;
assign io_out[1] = \io_out[1] ;
assign io_out[2] = \io_out[2] ;
assign io_out[3] = \io_out[3] ;
assign io_out[4] = \io_out[4] ;
assign io_out[5] = \io_out[5] ;
assign io_out[6] = \io_out[6] ;
assign io_out[7] = \io_out[7] ;
assign io_out[8] = \io_out[8] ;
assign io_out[9] = \io_out[9] ;
assign io_out[10] = \io_out[10] ;
assign io_out[11] = \io_out[11] ;
assign io_out[12] = \io_out[12] ;
assign io_out[13] = \io_out[13] ;
assign io_out[14] = \io_out[14] ;
assign io_out[15] = \io_out[15] ;
assign io_out[16] = \io_out[16] ;
assign io_out[17] = \io_out[17] ;
assign io_out[18] = \io_out[18] ;
assign io_out[19] = \io_out[19] ;
assign io_out[20] = \io_out[20] ;
assign io_out[21] = \io_out[21] ;
assign io_out[22] = \io_out[22] ;
assign io_out[23] = \io_out[23] ;
assign io_out[24] = \io_out[24] ;
assign io_out[25] = \io_out[25] ;
assign io_out[26] = \io_out[26] ;
assign io_out[27] = \io_out[27] ;
assign io_out[28] = \io_out[28] ;
assign io_out[29] = \io_out[29] ;
assign io_out[30] = \io_out[30] ;
assign io_out[31] = \io_out[31] ;
assign \io_sw[0] = io_sw[0] ;
assign \io_sw[1] = io_sw[1] ;
assign \io_sw[2] = io_sw[2] ;
assign \io_sw[3] = io_sw[3] ;

AND2_X1 _1811_ ( .A1(\io_in_b[31] ), .A2(fanout_net_1 ), .ZN(_0030_ ) );
NOR2_X1 _1812_ ( .A1(\io_in_b[31] ), .A2(fanout_net_1 ), .ZN(_0041_ ) );
NOR2_X1 _1813_ ( .A1(_0030_ ), .A2(_0041_ ), .ZN(_0052_ ) );
INV_X1 _1814_ ( .A(_0052_ ), .ZN(_0062_ ) );
XOR2_X1 _1815_ ( .A(\io_in_a[20] ), .B(\io_in_b[20] ), .Z(_0073_ ) );
XOR2_X2 _1816_ ( .A(\io_in_a[21] ), .B(\io_in_b[21] ), .Z(_0084_ ) );
NOR2_X1 _1817_ ( .A1(_0073_ ), .A2(_0084_ ), .ZN(_0095_ ) );
XOR2_X1 _1818_ ( .A(\io_in_b[23] ), .B(\io_in_a[23] ), .Z(_0105_ ) );
INV_X1 _1819_ ( .A(_0105_ ), .ZN(_0116_ ) );
XOR2_X1 _1820_ ( .A(\io_in_a[22] ), .B(\io_in_b[22] ), .Z(_0127_ ) );
INV_X1 _1821_ ( .A(_0127_ ), .ZN(_0138_ ) );
AND3_X1 _1822_ ( .A1(_0095_ ), .A2(_0116_ ), .A3(_0138_ ), .ZN(_0148_ ) );
XOR2_X1 _1823_ ( .A(\io_in_a[18] ), .B(\io_in_b[18] ), .Z(_0159_ ) );
AND2_X4 _1824_ ( .A1(\io_in_a[19] ), .A2(\io_in_b[19] ), .ZN(_0169_ ) );
NOR2_X1 _1825_ ( .A1(\io_in_a[19] ), .A2(\io_in_b[19] ), .ZN(_0180_ ) );
NOR2_X1 _1826_ ( .A1(_0169_ ), .A2(_0180_ ), .ZN(_0191_ ) );
NOR2_X1 _1827_ ( .A1(_0159_ ), .A2(_0191_ ), .ZN(_0202_ ) );
AND2_X4 _1828_ ( .A1(\io_in_a[17] ), .A2(\io_in_b[17] ), .ZN(_0213_ ) );
NOR2_X1 _1829_ ( .A1(\io_in_a[17] ), .A2(\io_in_b[17] ), .ZN(_0224_ ) );
NOR2_X4 _1830_ ( .A1(_0213_ ), .A2(_0224_ ), .ZN(_0234_ ) );
INV_X1 _1831_ ( .A(_0234_ ), .ZN(_0245_ ) );
AND2_X1 _1832_ ( .A1(\io_in_a[16] ), .A2(\io_in_b[16] ), .ZN(_0256_ ) );
NOR2_X1 _1833_ ( .A1(\io_in_a[16] ), .A2(\io_in_b[16] ), .ZN(_0267_ ) );
NOR2_X1 _1834_ ( .A1(_0256_ ), .A2(_0267_ ), .ZN(_0278_ ) );
INV_X1 _1835_ ( .A(_0278_ ), .ZN(_0289_ ) );
AND3_X1 _1836_ ( .A1(_0202_ ), .A2(_0245_ ), .A3(_0289_ ), .ZN(_0299_ ) );
AND2_X1 _1837_ ( .A1(_0148_ ), .A2(_0299_ ), .ZN(_0310_ ) );
INV_X1 _1838_ ( .A(_0310_ ), .ZN(_0321_ ) );
INV_X1 _1839_ ( .A(\io_in_a[7] ), .ZN(_0332_ ) );
NOR2_X1 _1840_ ( .A1(_0332_ ), .A2(\io_in_b[7] ), .ZN(_0342_ ) );
AND2_X4 _1841_ ( .A1(\io_in_b[5] ), .A2(\io_in_a[5] ), .ZN(_0353_ ) );
NOR2_X4 _1842_ ( .A1(\io_in_b[5] ), .A2(\io_in_a[5] ), .ZN(_0364_ ) );
NOR2_X4 _1843_ ( .A1(_0353_ ), .A2(_0364_ ), .ZN(_0374_ ) );
INV_X1 _1844_ ( .A(\io_in_a[4] ), .ZN(_0385_ ) );
NOR3_X4 _1845_ ( .A1(_0374_ ), .A2(\io_in_b[4] ), .A3(_0385_ ), .ZN(_0396_ ) );
INV_X1 _1846_ ( .A(\io_in_b[5] ), .ZN(_0406_ ) );
AOI21_X2 _1847_ ( .A(_0396_ ), .B1(_0406_ ), .B2(\io_in_a[5] ), .ZN(_0417_ ) );
XOR2_X1 _1848_ ( .A(\io_in_a[7] ), .B(\io_in_b[7] ), .Z(_0428_ ) );
XOR2_X1 _1849_ ( .A(\io_in_a[6] ), .B(\io_in_b[6] ), .Z(_0439_ ) );
NOR3_X1 _1850_ ( .A1(_0417_ ), .A2(_0428_ ), .A3(_0439_ ), .ZN(_0449_ ) );
INV_X1 _1851_ ( .A(_0428_ ), .ZN(_0460_ ) );
INV_X1 _1852_ ( .A(\io_in_a[6] ), .ZN(_0471_ ) );
NOR2_X1 _1853_ ( .A1(_0471_ ), .A2(\io_in_b[6] ), .ZN(_0482_ ) );
AOI211_X2 _1854_ ( .A(_0342_ ), .B(_0449_ ), .C1(_0460_ ), .C2(_0482_ ), .ZN(_0492_ ) );
INV_X1 _1855_ ( .A(\io_in_a[2] ), .ZN(_0503_ ) );
NOR2_X1 _1856_ ( .A1(_0503_ ), .A2(fanout_net_9 ), .ZN(_0514_ ) );
INV_X1 _1857_ ( .A(_0514_ ), .ZN(_0525_ ) );
INV_X1 _1858_ ( .A(\io_in_a[3] ), .ZN(_0535_ ) );
XOR2_X2 _1859_ ( .A(fanout_net_6 ), .B(\io_in_a[1] ), .Z(_0546_ ) );
INV_X1 _1860_ ( .A(fanout_net_3 ), .ZN(_0557_ ) );
NOR2_X1 _1861_ ( .A1(_0557_ ), .A2(\io_in_a[0] ), .ZN(_0567_ ) );
NOR2_X2 _1862_ ( .A1(_0546_ ), .A2(_0567_ ), .ZN(_0578_ ) );
INV_X1 _1863_ ( .A(fanout_net_6 ), .ZN(_0589_ ) );
AOI21_X2 _1864_ ( .A(_0578_ ), .B1(_0589_ ), .B2(\io_in_a[1] ), .ZN(_0600_ ) );
XOR2_X2 _1865_ ( .A(fanout_net_9 ), .B(\io_in_a[2] ), .Z(_0611_ ) );
OAI221_X1 _1866_ ( .A(_0525_ ), .B1(fanout_net_12 ), .B2(_0535_ ), .C1(_0600_ ), .C2(_0611_ ), .ZN(_0622_ ) );
NAND2_X1 _1867_ ( .A1(_0535_ ), .A2(fanout_net_12 ), .ZN(_0632_ ) );
XOR2_X1 _1868_ ( .A(\io_in_b[4] ), .B(\io_in_a[4] ), .Z(_0643_ ) );
NOR4_X1 _1869_ ( .A1(_0428_ ), .A2(_0439_ ), .A3(_0643_ ), .A4(_0374_ ), .ZN(_0654_ ) );
NAND3_X1 _1870_ ( .A1(_0622_ ), .A2(_0632_ ), .A3(_0654_ ), .ZN(_0664_ ) );
AND2_X2 _1871_ ( .A1(_0492_ ), .A2(_0664_ ), .ZN(_0675_ ) );
INV_X4 _1872_ ( .A(_0675_ ), .ZN(_0686_ ) );
XOR2_X1 _1873_ ( .A(\io_in_a[12] ), .B(\io_in_b[12] ), .Z(_0697_ ) );
AND2_X1 _1874_ ( .A1(\io_in_a[13] ), .A2(\io_in_b[13] ), .ZN(_0707_ ) );
NOR2_X1 _1875_ ( .A1(\io_in_a[13] ), .A2(\io_in_b[13] ), .ZN(_0718_ ) );
NOR2_X1 _1876_ ( .A1(_0707_ ), .A2(_0718_ ), .ZN(_0729_ ) );
NOR2_X1 _1877_ ( .A1(_0697_ ), .A2(_0729_ ), .ZN(_0739_ ) );
AND2_X1 _1878_ ( .A1(\io_in_a[15] ), .A2(\io_in_b[15] ), .ZN(_0750_ ) );
NOR2_X1 _1879_ ( .A1(\io_in_a[15] ), .A2(\io_in_b[15] ), .ZN(_0761_ ) );
NOR2_X1 _1880_ ( .A1(_0750_ ), .A2(_0761_ ), .ZN(_0771_ ) );
INV_X1 _1881_ ( .A(_0771_ ), .ZN(_0782_ ) );
XOR2_X1 _1882_ ( .A(\io_in_a[14] ), .B(\io_in_b[14] ), .Z(_0793_ ) );
INV_X1 _1883_ ( .A(_0793_ ), .ZN(_0803_ ) );
AND3_X1 _1884_ ( .A1(_0739_ ), .A2(_0782_ ), .A3(_0803_ ), .ZN(_0814_ ) );
XOR2_X1 _1885_ ( .A(\io_in_a[8] ), .B(\io_in_b[8] ), .Z(_0825_ ) );
AND2_X4 _1886_ ( .A1(\io_in_a[9] ), .A2(\io_in_b[9] ), .ZN(_0835_ ) );
NOR2_X4 _1887_ ( .A1(\io_in_a[9] ), .A2(\io_in_b[9] ), .ZN(_0846_ ) );
NOR2_X4 _1888_ ( .A1(_0835_ ), .A2(_0846_ ), .ZN(_0857_ ) );
NOR2_X1 _1889_ ( .A1(_0825_ ), .A2(_0857_ ), .ZN(_0867_ ) );
XOR2_X1 _1890_ ( .A(\io_in_a[10] ), .B(\io_in_b[10] ), .Z(_0878_ ) );
AND2_X4 _1891_ ( .A1(\io_in_a[11] ), .A2(\io_in_b[11] ), .ZN(_0889_ ) );
NOR2_X1 _1892_ ( .A1(\io_in_a[11] ), .A2(\io_in_b[11] ), .ZN(_0899_ ) );
NOR2_X1 _1893_ ( .A1(_0889_ ), .A2(_0899_ ), .ZN(_0910_ ) );
NOR2_X1 _1894_ ( .A1(_0878_ ), .A2(_0910_ ), .ZN(_0920_ ) );
NAND4_X4 _1895_ ( .A1(_0686_ ), .A2(_0814_ ), .A3(_0867_ ), .A4(_0920_ ), .ZN(_0931_ ) );
INV_X1 _1896_ ( .A(\io_in_a[8] ), .ZN(_0941_ ) );
NOR3_X4 _1897_ ( .A1(_0857_ ), .A2(_0941_ ), .A3(\io_in_b[8] ), .ZN(_0952_ ) );
INV_X1 _1898_ ( .A(\io_in_b[9] ), .ZN(_0963_ ) );
AOI21_X1 _1899_ ( .A(_0952_ ), .B1(\io_in_a[9] ), .B2(_0963_ ), .ZN(_0973_ ) );
NOR3_X1 _1900_ ( .A1(_0973_ ), .A2(_0910_ ), .A3(_0878_ ), .ZN(_0984_ ) );
INV_X1 _1901_ ( .A(\io_in_a[11] ), .ZN(_0994_ ) );
NOR2_X1 _1902_ ( .A1(_0994_ ), .A2(\io_in_b[11] ), .ZN(_1005_ ) );
INV_X1 _1903_ ( .A(\io_in_a[10] ), .ZN(_1012_ ) );
NOR3_X1 _1904_ ( .A1(_0910_ ), .A2(_1012_ ), .A3(\io_in_b[10] ), .ZN(_1013_ ) );
NOR3_X1 _1905_ ( .A1(_0984_ ), .A2(_1005_ ), .A3(_1013_ ), .ZN(_1014_ ) );
INV_X1 _1906_ ( .A(_1014_ ), .ZN(_1015_ ) );
NAND2_X1 _1907_ ( .A1(_1015_ ), .A2(_0814_ ), .ZN(_1016_ ) );
INV_X1 _1908_ ( .A(\io_in_a[12] ), .ZN(_1017_ ) );
NOR3_X1 _1909_ ( .A1(_0729_ ), .A2(_1017_ ), .A3(\io_in_b[12] ), .ZN(_1018_ ) );
INV_X1 _1910_ ( .A(\io_in_b[13] ), .ZN(_1019_ ) );
AOI21_X1 _1911_ ( .A(_1018_ ), .B1(\io_in_a[13] ), .B2(_1019_ ), .ZN(_1020_ ) );
OR3_X1 _1912_ ( .A1(_1020_ ), .A2(_0771_ ), .A3(_0793_ ), .ZN(_1021_ ) );
INV_X1 _1913_ ( .A(\io_in_a[15] ), .ZN(_1022_ ) );
OR2_X1 _1914_ ( .A1(_1022_ ), .A2(\io_in_b[15] ), .ZN(_1023_ ) );
INV_X1 _1915_ ( .A(\io_in_b[14] ), .ZN(_1024_ ) );
NAND3_X1 _1916_ ( .A1(_0782_ ), .A2(\io_in_a[14] ), .A3(_1024_ ), .ZN(_1025_ ) );
AND4_X4 _1917_ ( .A1(_1016_ ), .A2(_1021_ ), .A3(_1023_ ), .A4(_1025_ ), .ZN(_1026_ ) );
AOI21_X4 _1918_ ( .A(_0321_ ), .B1(_0931_ ), .B2(_1026_ ), .ZN(_1027_ ) );
INV_X1 _1919_ ( .A(\io_in_a[20] ), .ZN(_1028_ ) );
NOR3_X1 _1920_ ( .A1(_0084_ ), .A2(_1028_ ), .A3(\io_in_b[20] ), .ZN(_1029_ ) );
INV_X1 _1921_ ( .A(\io_in_b[21] ), .ZN(_1030_ ) );
AOI21_X1 _1922_ ( .A(_1029_ ), .B1(\io_in_a[21] ), .B2(_1030_ ), .ZN(_1031_ ) );
NOR3_X1 _1923_ ( .A1(_1031_ ), .A2(_0105_ ), .A3(_0127_ ), .ZN(_1032_ ) );
INV_X1 _1924_ ( .A(\io_in_a[22] ), .ZN(_1033_ ) );
NOR3_X1 _1925_ ( .A1(_0105_ ), .A2(_1033_ ), .A3(\io_in_b[22] ), .ZN(_1034_ ) );
INV_X1 _1926_ ( .A(\io_in_a[16] ), .ZN(_1035_ ) );
OR2_X1 _1927_ ( .A1(_1035_ ), .A2(\io_in_b[16] ), .ZN(_1036_ ) );
NOR2_X2 _1928_ ( .A1(_0234_ ), .A2(_1036_ ), .ZN(_1037_ ) );
INV_X1 _1929_ ( .A(\io_in_b[17] ), .ZN(_1038_ ) );
AOI21_X1 _1930_ ( .A(_1037_ ), .B1(\io_in_a[17] ), .B2(_1038_ ), .ZN(_1039_ ) );
NOR3_X1 _1931_ ( .A1(_1039_ ), .A2(_0191_ ), .A3(_0159_ ), .ZN(_1040_ ) );
INV_X1 _1932_ ( .A(\io_in_a[19] ), .ZN(_1041_ ) );
NOR2_X1 _1933_ ( .A1(_1041_ ), .A2(\io_in_b[19] ), .ZN(_1042_ ) );
INV_X1 _1934_ ( .A(\io_in_a[18] ), .ZN(_1043_ ) );
NOR3_X1 _1935_ ( .A1(_0191_ ), .A2(_1043_ ), .A3(\io_in_b[18] ), .ZN(_1044_ ) );
NOR3_X1 _1936_ ( .A1(_1040_ ), .A2(_1042_ ), .A3(_1044_ ), .ZN(_1045_ ) );
INV_X1 _1937_ ( .A(_1045_ ), .ZN(_1046_ ) );
AOI211_X1 _1938_ ( .A(_1032_ ), .B(_1034_ ), .C1(_1046_ ), .C2(_0148_ ), .ZN(_1047_ ) );
INV_X1 _1939_ ( .A(\io_in_a[23] ), .ZN(_1048_ ) );
OR2_X1 _1940_ ( .A1(_1048_ ), .A2(\io_in_b[23] ), .ZN(_1049_ ) );
AND2_X1 _1941_ ( .A1(_1047_ ), .A2(_1049_ ), .ZN(_1050_ ) );
INV_X2 _1942_ ( .A(_1050_ ), .ZN(_1051_ ) );
NOR2_X4 _1943_ ( .A1(_1027_ ), .A2(_1051_ ), .ZN(_1052_ ) );
XOR2_X1 _1944_ ( .A(\io_in_b[27] ), .B(\io_in_a[27] ), .Z(_1053_ ) );
INV_X1 _1945_ ( .A(_1053_ ), .ZN(_1054_ ) );
XOR2_X1 _1946_ ( .A(\io_in_b[26] ), .B(\io_in_a[26] ), .Z(_1055_ ) );
INV_X1 _1947_ ( .A(_1055_ ), .ZN(_1056_ ) );
NAND2_X1 _1948_ ( .A1(_1054_ ), .A2(_1056_ ), .ZN(_1057_ ) );
AND2_X1 _1949_ ( .A1(\io_in_b[25] ), .A2(\io_in_a[25] ), .ZN(_1058_ ) );
NOR2_X1 _1950_ ( .A1(\io_in_b[25] ), .A2(\io_in_a[25] ), .ZN(_1059_ ) );
NOR2_X1 _1951_ ( .A1(_1058_ ), .A2(_1059_ ), .ZN(_1060_ ) );
XOR2_X1 _1952_ ( .A(\io_in_b[24] ), .B(\io_in_a[24] ), .Z(_1061_ ) );
NOR4_X2 _1953_ ( .A1(_1052_ ), .A2(_1057_ ), .A3(_1060_ ), .A4(_1061_ ), .ZN(_1062_ ) );
INV_X1 _1954_ ( .A(\io_in_a[27] ), .ZN(_1063_ ) );
NOR2_X1 _1955_ ( .A1(_1063_ ), .A2(\io_in_b[27] ), .ZN(_1064_ ) );
INV_X1 _1956_ ( .A(\io_in_a[26] ), .ZN(_1065_ ) );
OR3_X1 _1957_ ( .A1(_1053_ ), .A2(\io_in_b[26] ), .A3(_1065_ ), .ZN(_1066_ ) );
INV_X1 _1958_ ( .A(\io_in_a[24] ), .ZN(_1067_ ) );
NOR3_X1 _1959_ ( .A1(_1060_ ), .A2(\io_in_b[24] ), .A3(_1067_ ), .ZN(_1068_ ) );
INV_X1 _1960_ ( .A(\io_in_a[25] ), .ZN(_1069_ ) );
NOR2_X1 _1961_ ( .A1(_1069_ ), .A2(\io_in_b[25] ), .ZN(_1070_ ) );
NOR2_X1 _1962_ ( .A1(_1068_ ), .A2(_1070_ ), .ZN(_1071_ ) );
OAI21_X1 _1963_ ( .A(_1066_ ), .B1(_1071_ ), .B2(_1057_ ), .ZN(_1072_ ) );
OR3_X4 _1964_ ( .A1(_1062_ ), .A2(_1064_ ), .A3(_1072_ ), .ZN(_1073_ ) );
XOR2_X1 _1965_ ( .A(\io_in_a[30] ), .B(\io_in_b[30] ), .Z(_1074_ ) );
INV_X1 _1966_ ( .A(_1074_ ), .ZN(_1075_ ) );
XOR2_X1 _1967_ ( .A(\io_in_b[28] ), .B(\io_in_a[28] ), .Z(_1076_ ) );
AND2_X1 _1968_ ( .A1(\io_in_b[29] ), .A2(\io_in_a[29] ), .ZN(_1077_ ) );
NOR2_X1 _1969_ ( .A1(\io_in_b[29] ), .A2(\io_in_a[29] ), .ZN(_1078_ ) );
NOR2_X1 _1970_ ( .A1(_1077_ ), .A2(_1078_ ), .ZN(_1079_ ) );
NOR2_X1 _1971_ ( .A1(_1076_ ), .A2(_1079_ ), .ZN(_1080_ ) );
AND4_X4 _1972_ ( .A1(_0062_ ), .A2(_1073_ ), .A3(_1075_ ), .A4(_1080_ ), .ZN(_1081_ ) );
INV_X1 _1973_ ( .A(fanout_net_1 ), .ZN(_1082_ ) );
NOR2_X1 _1974_ ( .A1(_1082_ ), .A2(\io_in_b[31] ), .ZN(_1083_ ) );
INV_X1 _1975_ ( .A(\io_in_a[28] ), .ZN(_1084_ ) );
NOR3_X1 _1976_ ( .A1(_1079_ ), .A2(\io_in_b[28] ), .A3(_1084_ ), .ZN(_1085_ ) );
INV_X1 _1977_ ( .A(_1085_ ), .ZN(_1086_ ) );
INV_X1 _1978_ ( .A(\io_in_a[29] ), .ZN(_1087_ ) );
OAI21_X1 _1979_ ( .A(_1086_ ), .B1(\io_in_b[29] ), .B2(_1087_ ), .ZN(_1088_ ) );
AND3_X1 _1980_ ( .A1(_1088_ ), .A2(_0062_ ), .A3(_1075_ ), .ZN(_1089_ ) );
OR3_X4 _1981_ ( .A1(_1081_ ), .A2(_1083_ ), .A3(_1089_ ), .ZN(_1090_ ) );
INV_X1 _1982_ ( .A(\io_in_a[30] ), .ZN(_1091_ ) );
NOR3_X1 _1983_ ( .A1(_0052_ ), .A2(_1091_ ), .A3(\io_in_b[30] ), .ZN(_1092_ ) );
INV_X1 _1984_ ( .A(\io_sw[3] ), .ZN(_1093_ ) );
INV_X1 _1985_ ( .A(\io_sw[2] ), .ZN(_1094_ ) );
INV_X1 _1986_ ( .A(\io_sw[1] ), .ZN(_1095_ ) );
NAND3_X1 _1987_ ( .A1(_1093_ ), .A2(_1094_ ), .A3(_1095_ ), .ZN(_1096_ ) );
INV_X1 _1988_ ( .A(\io_sw[0] ), .ZN(_1097_ ) );
NOR2_X1 _1989_ ( .A1(_1096_ ), .A2(_1097_ ), .ZN(_1098_ ) );
INV_X1 _1990_ ( .A(_1098_ ), .ZN(_1099_ ) );
BUF_X2 _1991_ ( .A(_1099_ ), .Z(_1100_ ) );
BUF_X2 _1992_ ( .A(_1100_ ), .Z(_1101_ ) );
OR3_X1 _1993_ ( .A1(_1090_ ), .A2(_1092_ ), .A3(_1101_ ), .ZN(_1102_ ) );
NOR2_X1 _1994_ ( .A1(\io_sw[3] ), .A2(\io_sw[2] ), .ZN(_1103_ ) );
NOR2_X1 _1995_ ( .A1(\io_sw[0] ), .A2(\io_sw[1] ), .ZN(_1104_ ) );
AND2_X2 _1996_ ( .A1(_1103_ ), .A2(_1104_ ), .ZN(_1105_ ) );
BUF_X2 _1997_ ( .A(_1105_ ), .Z(_1106_ ) );
INV_X1 _1998_ ( .A(_1059_ ), .ZN(_1107_ ) );
AND2_X1 _1999_ ( .A1(\io_in_b[24] ), .A2(\io_in_a[24] ), .ZN(_1108_ ) );
AOI21_X1 _2000_ ( .A(_1058_ ), .B1(_1107_ ), .B2(_1108_ ), .ZN(_1109_ ) );
OR3_X1 _2001_ ( .A1(_1054_ ), .A2(_1056_ ), .A3(_1109_ ), .ZN(_1110_ ) );
AND2_X1 _2002_ ( .A1(\io_in_b[27] ), .A2(\io_in_a[27] ), .ZN(_1111_ ) );
AND2_X1 _2003_ ( .A1(\io_in_b[26] ), .A2(\io_in_a[26] ), .ZN(_1112_ ) );
AOI21_X1 _2004_ ( .A(_1111_ ), .B1(_1053_ ), .B2(_1112_ ), .ZN(_1113_ ) );
NAND2_X1 _2005_ ( .A1(_1110_ ), .A2(_1113_ ), .ZN(_1114_ ) );
AND2_X1 _2006_ ( .A1(\io_in_a[7] ), .A2(\io_in_b[7] ), .ZN(_1115_ ) );
INV_X1 _2007_ ( .A(_0439_ ), .ZN(_1116_ ) );
AND2_X1 _2008_ ( .A1(\io_in_b[4] ), .A2(\io_in_a[4] ), .ZN(_1117_ ) );
NOR2_X1 _2009_ ( .A1(_1117_ ), .A2(_0353_ ), .ZN(_1118_ ) );
NOR4_X1 _2010_ ( .A1(_0460_ ), .A2(_1116_ ), .A3(_0364_ ), .A4(_1118_ ), .ZN(_1119_ ) );
AND2_X1 _2011_ ( .A1(\io_in_a[6] ), .A2(\io_in_b[6] ), .ZN(_1120_ ) );
AOI211_X1 _2012_ ( .A(_1115_ ), .B(_1119_ ), .C1(_0428_ ), .C2(_1120_ ), .ZN(_1121_ ) );
AND2_X1 _2013_ ( .A1(fanout_net_6 ), .A2(\io_in_a[1] ), .ZN(_1122_ ) );
AND2_X1 _2014_ ( .A1(\io_in_a[0] ), .A2(fanout_net_3 ), .ZN(_1123_ ) );
AOI21_X4 _2015_ ( .A(_1122_ ), .B1(_0546_ ), .B2(_1123_ ), .ZN(_1124_ ) );
INV_X1 _2016_ ( .A(_0611_ ), .ZN(_1125_ ) );
AND2_X4 _2017_ ( .A1(fanout_net_12 ), .A2(\io_in_a[3] ), .ZN(_1126_ ) );
NOR2_X1 _2018_ ( .A1(fanout_net_12 ), .A2(\io_in_a[3] ), .ZN(_1127_ ) );
NOR2_X1 _2019_ ( .A1(_1126_ ), .A2(_1127_ ), .ZN(_1128_ ) );
INV_X1 _2020_ ( .A(_1128_ ), .ZN(_1129_ ) );
OR3_X2 _2021_ ( .A1(_1124_ ), .A2(_1125_ ), .A3(_1129_ ), .ZN(_1130_ ) );
AND2_X1 _2022_ ( .A1(fanout_net_9 ), .A2(\io_in_a[2] ), .ZN(_1131_ ) );
AOI21_X1 _2023_ ( .A(_1126_ ), .B1(_1128_ ), .B2(_1131_ ), .ZN(_1132_ ) );
NAND2_X2 _2024_ ( .A1(_1130_ ), .A2(_1132_ ), .ZN(_1133_ ) );
AND4_X1 _2025_ ( .A1(_0428_ ), .A2(_0439_ ), .A3(_0643_ ), .A4(_0374_ ), .ZN(_1134_ ) );
NAND2_X1 _2026_ ( .A1(_1133_ ), .A2(_1134_ ), .ZN(_1135_ ) );
NAND2_X2 _2027_ ( .A1(_1121_ ), .A2(_1135_ ), .ZN(_1136_ ) );
AND2_X1 _2028_ ( .A1(_0793_ ), .A2(_0771_ ), .ZN(_1137_ ) );
AND2_X1 _2029_ ( .A1(_0697_ ), .A2(_0729_ ), .ZN(_1138_ ) );
AND2_X1 _2030_ ( .A1(_1137_ ), .A2(_1138_ ), .ZN(_1139_ ) );
AND2_X1 _2031_ ( .A1(_0825_ ), .A2(_0857_ ), .ZN(_1140_ ) );
AND2_X1 _2032_ ( .A1(_0878_ ), .A2(_0910_ ), .ZN(_1141_ ) );
NAND4_X1 _2033_ ( .A1(_1136_ ), .A2(_1139_ ), .A3(_1140_ ), .A4(_1141_ ), .ZN(_1142_ ) );
INV_X1 _2034_ ( .A(_1139_ ), .ZN(_1143_ ) );
AND2_X1 _2035_ ( .A1(\io_in_a[8] ), .A2(\io_in_b[8] ), .ZN(_1144_ ) );
AOI21_X1 _2036_ ( .A(_0835_ ), .B1(_0857_ ), .B2(_1144_ ), .ZN(_1145_ ) );
INV_X1 _2037_ ( .A(_1145_ ), .ZN(_1146_ ) );
NAND2_X1 _2038_ ( .A1(_1146_ ), .A2(_1141_ ), .ZN(_1147_ ) );
INV_X1 _2039_ ( .A(_0889_ ), .ZN(_1148_ ) );
AND2_X1 _2040_ ( .A1(\io_in_a[10] ), .A2(\io_in_b[10] ), .ZN(_1149_ ) );
INV_X1 _2041_ ( .A(_1149_ ), .ZN(_1150_ ) );
AOI21_X1 _2042_ ( .A(_0899_ ), .B1(_1148_ ), .B2(_1150_ ), .ZN(_1151_ ) );
INV_X1 _2043_ ( .A(_1151_ ), .ZN(_1152_ ) );
AOI21_X1 _2044_ ( .A(_1143_ ), .B1(_1147_ ), .B2(_1152_ ), .ZN(_1153_ ) );
AND2_X1 _2045_ ( .A1(\io_in_a[12] ), .A2(\io_in_b[12] ), .ZN(_1154_ ) );
AOI21_X1 _2046_ ( .A(_0707_ ), .B1(_0729_ ), .B2(_1154_ ), .ZN(_1155_ ) );
NOR3_X1 _2047_ ( .A1(_1155_ ), .A2(_0803_ ), .A3(_0782_ ), .ZN(_1156_ ) );
AND2_X1 _2048_ ( .A1(\io_in_a[14] ), .A2(\io_in_b[14] ), .ZN(_1157_ ) );
INV_X1 _2049_ ( .A(_1157_ ), .ZN(_1158_ ) );
NOR3_X1 _2050_ ( .A1(_1158_ ), .A2(_0750_ ), .A3(_0761_ ), .ZN(_1159_ ) );
NOR4_X1 _2051_ ( .A1(_1153_ ), .A2(_0750_ ), .A3(_1156_ ), .A4(_1159_ ), .ZN(_1160_ ) );
AND2_X2 _2052_ ( .A1(_1142_ ), .A2(_1160_ ), .ZN(_1161_ ) );
INV_X2 _2053_ ( .A(_1161_ ), .ZN(_1162_ ) );
AND2_X1 _2054_ ( .A1(_0073_ ), .A2(_0084_ ), .ZN(_1163_ ) );
AND3_X1 _2055_ ( .A1(_1163_ ), .A2(_0105_ ), .A3(_0127_ ), .ZN(_1164_ ) );
AND2_X1 _2056_ ( .A1(_0159_ ), .A2(_0191_ ), .ZN(_1165_ ) );
AND2_X1 _2057_ ( .A1(_0234_ ), .A2(_0278_ ), .ZN(_1166_ ) );
NAND4_X4 _2058_ ( .A1(_1162_ ), .A2(_1164_ ), .A3(_1165_ ), .A4(_1166_ ), .ZN(_1167_ ) );
INV_X1 _2059_ ( .A(_0180_ ), .ZN(_1168_ ) );
AND2_X1 _2060_ ( .A1(\io_in_a[18] ), .A2(\io_in_b[18] ), .ZN(_1169_ ) );
OAI21_X1 _2061_ ( .A(_1168_ ), .B1(_0169_ ), .B2(_1169_ ), .ZN(_1170_ ) );
INV_X1 _2062_ ( .A(_1165_ ), .ZN(_1171_ ) );
AOI21_X1 _2063_ ( .A(_0213_ ), .B1(_0234_ ), .B2(_0256_ ), .ZN(_1172_ ) );
OAI21_X1 _2064_ ( .A(_1170_ ), .B1(_1171_ ), .B2(_1172_ ), .ZN(_1173_ ) );
NAND2_X1 _2065_ ( .A1(_1173_ ), .A2(_1164_ ), .ZN(_1174_ ) );
AND2_X1 _2066_ ( .A1(\io_in_a[21] ), .A2(\io_in_b[21] ), .ZN(_1175_ ) );
AND2_X1 _2067_ ( .A1(\io_in_a[20] ), .A2(\io_in_b[20] ), .ZN(_1176_ ) );
AOI21_X1 _2068_ ( .A(_1175_ ), .B1(_0084_ ), .B2(_1176_ ), .ZN(_1177_ ) );
OR3_X1 _2069_ ( .A1(_1177_ ), .A2(_0116_ ), .A3(_0138_ ), .ZN(_1178_ ) );
AND2_X1 _2070_ ( .A1(\io_in_b[23] ), .A2(\io_in_a[23] ), .ZN(_1179_ ) );
AND2_X1 _2071_ ( .A1(\io_in_a[22] ), .A2(\io_in_b[22] ), .ZN(_1180_ ) );
AOI21_X1 _2072_ ( .A(_1179_ ), .B1(_0105_ ), .B2(_1180_ ), .ZN(_1181_ ) );
AND3_X1 _2073_ ( .A1(_1174_ ), .A2(_1178_ ), .A3(_1181_ ), .ZN(_1182_ ) );
NAND2_X1 _2074_ ( .A1(_1167_ ), .A2(_1182_ ), .ZN(_1183_ ) );
AND2_X1 _2075_ ( .A1(_1061_ ), .A2(_1060_ ), .ZN(_1184_ ) );
AND3_X1 _2076_ ( .A1(_1184_ ), .A2(_1053_ ), .A3(_1055_ ), .ZN(_1185_ ) );
AOI21_X2 _2077_ ( .A(_1114_ ), .B1(_1183_ ), .B2(_1185_ ), .ZN(_1186_ ) );
INV_X1 _2078_ ( .A(_1079_ ), .ZN(_1187_ ) );
INV_X1 _2079_ ( .A(_1076_ ), .ZN(_1188_ ) );
OR3_X4 _2080_ ( .A1(_1186_ ), .A2(_1187_ ), .A3(_1188_ ), .ZN(_1189_ ) );
NAND2_X1 _2081_ ( .A1(_1074_ ), .A2(_0052_ ), .ZN(_1190_ ) );
NOR2_X1 _2082_ ( .A1(_1189_ ), .A2(_1190_ ), .ZN(_1191_ ) );
AND2_X1 _2083_ ( .A1(\io_in_b[28] ), .A2(\io_in_a[28] ), .ZN(_1192_ ) );
AOI21_X1 _2084_ ( .A(_1077_ ), .B1(_1079_ ), .B2(_1192_ ), .ZN(_1193_ ) );
NOR2_X1 _2085_ ( .A1(_1193_ ), .A2(_1190_ ), .ZN(_1194_ ) );
AND2_X1 _2086_ ( .A1(\io_in_a[30] ), .A2(\io_in_b[30] ), .ZN(_1195_ ) );
INV_X1 _2087_ ( .A(_1195_ ), .ZN(_1196_ ) );
NOR2_X1 _2088_ ( .A1(_1196_ ), .A2(_0041_ ), .ZN(_1197_ ) );
OR3_X1 _2089_ ( .A1(_1194_ ), .A2(_0030_ ), .A3(_1197_ ), .ZN(_1198_ ) );
OAI21_X1 _2090_ ( .A(_1106_ ), .B1(_1191_ ), .B2(_1198_ ), .ZN(_1199_ ) );
NAND2_X1 _2091_ ( .A1(_1102_ ), .A2(_1199_ ), .ZN(io_carry ) );
NAND4_X1 _2092_ ( .A1(_1093_ ), .A2(_1094_ ), .A3(_1097_ ), .A4(\io_sw[1] ), .ZN(_1200_ ) );
NOR3_X1 _2093_ ( .A1(_1090_ ), .A2(_1092_ ), .A3(_1200_ ), .ZN(_1201_ ) );
INV_X1 _2094_ ( .A(\io_in_b[4] ), .ZN(_1202_ ) );
BUF_X4 _2095_ ( .A(_1202_ ), .Z(_1203_ ) );
BUF_X4 _2096_ ( .A(_0557_ ), .Z(_1204_ ) );
BUF_X4 _2097_ ( .A(_1204_ ), .Z(_1205_ ) );
BUF_X2 _2098_ ( .A(_1205_ ), .Z(_1206_ ) );
AND2_X1 _2099_ ( .A1(_1206_ ), .A2(\io_in_a[0] ), .ZN(_1207_ ) );
INV_X2 _2100_ ( .A(fanout_net_9 ), .ZN(_1208_ ) );
BUF_X4 _2101_ ( .A(_1208_ ), .Z(_1209_ ) );
BUF_X4 _2102_ ( .A(_0589_ ), .Z(_1210_ ) );
BUF_X4 _2103_ ( .A(_1210_ ), .Z(_1211_ ) );
BUF_X2 _2104_ ( .A(_1211_ ), .Z(_1212_ ) );
AND3_X1 _2105_ ( .A1(_1207_ ), .A2(_1209_ ), .A3(_1212_ ), .ZN(_1213_ ) );
INV_X2 _2106_ ( .A(fanout_net_12 ), .ZN(_1214_ ) );
BUF_X4 _2107_ ( .A(_1214_ ), .Z(_1215_ ) );
BUF_X2 _2108_ ( .A(_1215_ ), .Z(_1216_ ) );
NOR2_X1 _2109_ ( .A1(_1093_ ), .A2(\io_sw[2] ), .ZN(_1217_ ) );
AND2_X1 _2110_ ( .A1(_1217_ ), .A2(_1104_ ), .ZN(_1218_ ) );
AND4_X1 _2111_ ( .A1(_1203_ ), .A2(_1213_ ), .A3(_1216_ ), .A4(_1218_ ), .ZN(_1219_ ) );
NOR2_X1 _2112_ ( .A1(\io_in_a[0] ), .A2(fanout_net_3 ), .ZN(_1220_ ) );
NOR2_X1 _2113_ ( .A1(_1094_ ), .A2(\io_sw[3] ), .ZN(_1221_ ) );
BUF_X2 _2114_ ( .A(_1221_ ), .Z(_1222_ ) );
AND2_X2 _2115_ ( .A1(_1222_ ), .A2(_1104_ ), .ZN(_1223_ ) );
INV_X1 _2116_ ( .A(_1223_ ), .ZN(_1224_ ) );
AOI211_X1 _2117_ ( .A(_1123_ ), .B(_1220_ ), .C1(_1224_ ), .C2(_1096_ ), .ZN(_1225_ ) );
NOR2_X1 _2118_ ( .A1(_1095_ ), .A2(\io_sw[0] ), .ZN(_1226_ ) );
AND2_X1 _2119_ ( .A1(_1226_ ), .A2(_1222_ ), .ZN(_1227_ ) );
BUF_X4 _2120_ ( .A(_1227_ ), .Z(_1228_ ) );
INV_X1 _2121_ ( .A(_1228_ ), .ZN(_1229_ ) );
INV_X1 _2122_ ( .A(_1123_ ), .ZN(_1230_ ) );
AND2_X1 _2123_ ( .A1(\io_sw[0] ), .A2(\io_sw[1] ), .ZN(_1231_ ) );
AND2_X1 _2124_ ( .A1(_1231_ ), .A2(_1103_ ), .ZN(_1232_ ) );
INV_X1 _2125_ ( .A(_1232_ ), .ZN(_1233_ ) );
BUF_X4 _2126_ ( .A(_1233_ ), .Z(_1234_ ) );
OAI22_X1 _2127_ ( .A1(_1229_ ), .A2(_1230_ ), .B1(_1234_ ), .B2(_1220_ ), .ZN(_1235_ ) );
NOR4_X1 _2128_ ( .A1(_1201_ ), .A2(_1219_ ), .A3(_1225_ ), .A4(_1235_ ), .ZN(_1236_ ) );
NOR2_X1 _2129_ ( .A1(_1097_ ), .A2(\io_sw[1] ), .ZN(_1237_ ) );
AND2_X2 _2130_ ( .A1(_1237_ ), .A2(_1217_ ), .ZN(_1238_ ) );
AND2_X1 _2131_ ( .A1(_1238_ ), .A2(_0406_ ), .ZN(_1239_ ) );
BUF_X4 _2132_ ( .A(_1210_ ), .Z(_1240_ ) );
NOR2_X1 _2133_ ( .A1(\io_in_b[31] ), .A2(\io_in_b[29] ), .ZN(_1241_ ) );
INV_X1 _2134_ ( .A(\io_in_b[12] ), .ZN(_1242_ ) );
AND3_X1 _2135_ ( .A1(_1241_ ), .A2(_1019_ ), .A3(_1242_ ), .ZN(_1243_ ) );
NAND3_X1 _2136_ ( .A1(_1243_ ), .A2(_1038_ ), .A3(_1024_ ), .ZN(_1244_ ) );
OR2_X4 _2137_ ( .A1(\io_in_b[24] ), .A2(\io_in_b[23] ), .ZN(_1245_ ) );
OR3_X4 _2138_ ( .A1(_1245_ ), .A2(\io_in_b[11] ), .A3(\io_in_b[10] ), .ZN(_1246_ ) );
NOR4_X4 _2139_ ( .A1(_1244_ ), .A2(_1246_ ), .A3(\io_in_b[28] ), .A4(\io_in_b[25] ), .ZN(_1247_ ) );
NOR4_X1 _2140_ ( .A1(\io_in_b[30] ), .A2(\io_in_b[22] ), .A3(\io_in_b[21] ), .A4(\io_in_b[18] ), .ZN(_1248_ ) );
NOR4_X1 _2141_ ( .A1(\io_in_b[20] ), .A2(\io_in_b[19] ), .A3(\io_in_b[16] ), .A4(\io_in_b[15] ), .ZN(_1249_ ) );
NAND2_X1 _2142_ ( .A1(_1248_ ), .A2(_1249_ ), .ZN(_1250_ ) );
OR2_X4 _2143_ ( .A1(\io_in_b[9] ), .A2(\io_in_b[6] ), .ZN(_1251_ ) );
OR3_X4 _2144_ ( .A1(_1251_ ), .A2(\io_in_b[8] ), .A3(\io_in_b[7] ), .ZN(_1252_ ) );
NOR4_X4 _2145_ ( .A1(_1250_ ), .A2(_1252_ ), .A3(\io_in_b[27] ), .A4(\io_in_b[26] ), .ZN(_1253_ ) );
AND2_X2 _2146_ ( .A1(_1247_ ), .A2(_1253_ ), .ZN(_1254_ ) );
BUF_X4 _2147_ ( .A(_1254_ ), .Z(_1255_ ) );
INV_X1 _2148_ ( .A(_1255_ ), .ZN(_1256_ ) );
BUF_X4 _2149_ ( .A(_1256_ ), .Z(_1257_ ) );
NAND2_X1 _2150_ ( .A1(fanout_net_3 ), .A2(\io_in_a[27] ), .ZN(_1258_ ) );
BUF_X4 _2151_ ( .A(_1205_ ), .Z(_1259_ ) );
NAND2_X1 _2152_ ( .A1(_1259_ ), .A2(\io_in_a[26] ), .ZN(_1260_ ) );
AOI211_X1 _2153_ ( .A(_1240_ ), .B(_1257_ ), .C1(_1258_ ), .C2(_1260_ ), .ZN(_1261_ ) );
INV_X1 _2154_ ( .A(_1261_ ), .ZN(_1262_ ) );
NAND2_X1 _2155_ ( .A1(fanout_net_3 ), .A2(\io_in_a[25] ), .ZN(_1263_ ) );
NOR2_X1 _2156_ ( .A1(_1067_ ), .A2(fanout_net_3 ), .ZN(_1264_ ) );
INV_X1 _2157_ ( .A(_1264_ ), .ZN(_1265_ ) );
AOI211_X1 _2158_ ( .A(fanout_net_6 ), .B(_1257_ ), .C1(_1263_ ), .C2(_1265_ ), .ZN(_1266_ ) );
INV_X1 _2159_ ( .A(_1266_ ), .ZN(_1267_ ) );
AOI21_X1 _2160_ ( .A(fanout_net_9 ), .B1(_1262_ ), .B2(_1267_ ), .ZN(_1268_ ) );
BUF_X4 _2161_ ( .A(_1255_ ), .Z(_1269_ ) );
AND2_X1 _2162_ ( .A1(fanout_net_3 ), .A2(fanout_net_1 ), .ZN(_1270_ ) );
NOR2_X1 _2163_ ( .A1(_1091_ ), .A2(fanout_net_3 ), .ZN(_1271_ ) );
OAI21_X1 _2164_ ( .A(_1269_ ), .B1(_1270_ ), .B2(_1271_ ), .ZN(_1272_ ) );
NOR2_X1 _2165_ ( .A1(_1272_ ), .A2(_1240_ ), .ZN(_1273_ ) );
NAND2_X1 _2166_ ( .A1(fanout_net_3 ), .A2(\io_in_a[29] ), .ZN(_1274_ ) );
BUF_X4 _2167_ ( .A(_1204_ ), .Z(_1275_ ) );
NAND2_X1 _2168_ ( .A1(_1275_ ), .A2(\io_in_a[28] ), .ZN(_1276_ ) );
AOI21_X1 _2169_ ( .A(_1257_ ), .B1(_1274_ ), .B2(_1276_ ), .ZN(_1277_ ) );
AOI21_X1 _2170_ ( .A(_1273_ ), .B1(_1212_ ), .B2(_1277_ ), .ZN(_1278_ ) );
BUF_X4 _2171_ ( .A(_1209_ ), .Z(_1279_ ) );
NOR2_X1 _2172_ ( .A1(_1278_ ), .A2(_1279_ ), .ZN(_1280_ ) );
OAI21_X1 _2173_ ( .A(fanout_net_12 ), .B1(_1268_ ), .B2(_1280_ ), .ZN(_1281_ ) );
BUF_X4 _2174_ ( .A(_1214_ ), .Z(_1282_ ) );
BUF_X4 _2175_ ( .A(_1282_ ), .Z(_1283_ ) );
BUF_X4 _2176_ ( .A(_1209_ ), .Z(_1284_ ) );
BUF_X4 _2177_ ( .A(_1255_ ), .Z(_1285_ ) );
BUF_X4 _2178_ ( .A(_1285_ ), .Z(_1286_ ) );
NOR2_X1 _2179_ ( .A1(_1033_ ), .A2(fanout_net_3 ), .ZN(_1287_ ) );
AND2_X1 _2180_ ( .A1(fanout_net_3 ), .A2(\io_in_a[23] ), .ZN(_1288_ ) );
OAI211_X1 _2181_ ( .A(_1286_ ), .B(fanout_net_6 ), .C1(_1287_ ), .C2(_1288_ ), .ZN(_1289_ ) );
BUF_X4 _2182_ ( .A(_0589_ ), .Z(_1290_ ) );
BUF_X4 _2183_ ( .A(_1290_ ), .Z(_1291_ ) );
AND2_X1 _2184_ ( .A1(fanout_net_3 ), .A2(\io_in_a[21] ), .ZN(_1292_ ) );
NOR2_X1 _2185_ ( .A1(_1028_ ), .A2(fanout_net_3 ), .ZN(_1293_ ) );
OAI211_X1 _2186_ ( .A(_1286_ ), .B(_1291_ ), .C1(_1292_ ), .C2(_1293_ ), .ZN(_1294_ ) );
AOI21_X1 _2187_ ( .A(_1284_ ), .B1(_1289_ ), .B2(_1294_ ), .ZN(_1295_ ) );
BUF_X8 _2188_ ( .A(_1255_ ), .Z(_1296_ ) );
BUF_X4 _2189_ ( .A(_1296_ ), .Z(_1297_ ) );
BUF_X4 _2190_ ( .A(_1297_ ), .Z(_1298_ ) );
AND2_X1 _2191_ ( .A1(fanout_net_3 ), .A2(\io_in_a[19] ), .ZN(_1299_ ) );
NOR2_X1 _2192_ ( .A1(_1043_ ), .A2(fanout_net_3 ), .ZN(_1300_ ) );
OAI211_X1 _2193_ ( .A(_1298_ ), .B(fanout_net_6 ), .C1(_1299_ ), .C2(_1300_ ), .ZN(_1301_ ) );
AND2_X1 _2194_ ( .A1(fanout_net_3 ), .A2(\io_in_a[17] ), .ZN(_1302_ ) );
NOR2_X1 _2195_ ( .A1(_1035_ ), .A2(fanout_net_3 ), .ZN(_1303_ ) );
OAI211_X1 _2196_ ( .A(_1298_ ), .B(_1212_ ), .C1(_1302_ ), .C2(_1303_ ), .ZN(_1304_ ) );
AOI21_X1 _2197_ ( .A(fanout_net_9 ), .B1(_1301_ ), .B2(_1304_ ), .ZN(_1305_ ) );
OAI21_X1 _2198_ ( .A(_1283_ ), .B1(_1295_ ), .B2(_1305_ ), .ZN(_1306_ ) );
NAND2_X1 _2199_ ( .A1(_1281_ ), .A2(_1306_ ), .ZN(_1307_ ) );
BUF_X4 _2200_ ( .A(_1247_ ), .Z(_1308_ ) );
BUF_X4 _2201_ ( .A(_1308_ ), .Z(_1309_ ) );
BUF_X2 _2202_ ( .A(_1309_ ), .Z(_1310_ ) );
BUF_X4 _2203_ ( .A(_1253_ ), .Z(_1311_ ) );
BUF_X4 _2204_ ( .A(_1311_ ), .Z(_1312_ ) );
BUF_X2 _2205_ ( .A(_1312_ ), .Z(_1313_ ) );
MUX2_X1 _2206_ ( .A(\io_in_a[8] ), .B(\io_in_a[9] ), .S(fanout_net_3 ), .Z(_1314_ ) );
NAND4_X1 _2207_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1240_ ), .A4(_1314_ ), .ZN(_1315_ ) );
MUX2_X1 _2208_ ( .A(\io_in_a[10] ), .B(\io_in_a[11] ), .S(fanout_net_3 ), .Z(_1316_ ) );
NAND3_X1 _2209_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1316_ ), .ZN(_1317_ ) );
BUF_X4 _2210_ ( .A(_1211_ ), .Z(_1318_ ) );
OAI21_X1 _2211_ ( .A(_1315_ ), .B1(_1317_ ), .B2(_1318_ ), .ZN(_1319_ ) );
BUF_X4 _2212_ ( .A(_1208_ ), .Z(_1320_ ) );
BUF_X4 _2213_ ( .A(_1320_ ), .Z(_1321_ ) );
NAND2_X1 _2214_ ( .A1(_1319_ ), .A2(_1321_ ), .ZN(_1322_ ) );
AND2_X1 _2215_ ( .A1(fanout_net_3 ), .A2(\io_in_a[15] ), .ZN(_1323_ ) );
INV_X1 _2216_ ( .A(\io_in_a[14] ), .ZN(_1324_ ) );
NOR2_X1 _2217_ ( .A1(_1324_ ), .A2(fanout_net_3 ), .ZN(_1325_ ) );
OAI211_X1 _2218_ ( .A(_1286_ ), .B(fanout_net_6 ), .C1(_1323_ ), .C2(_1325_ ), .ZN(_1326_ ) );
BUF_X4 _2219_ ( .A(_1290_ ), .Z(_1327_ ) );
AND2_X1 _2220_ ( .A1(fanout_net_3 ), .A2(\io_in_a[13] ), .ZN(_1328_ ) );
NOR2_X1 _2221_ ( .A1(_1017_ ), .A2(fanout_net_3 ), .ZN(_1329_ ) );
OAI211_X1 _2222_ ( .A(_1286_ ), .B(_1327_ ), .C1(_1328_ ), .C2(_1329_ ), .ZN(_1330_ ) );
AND2_X1 _2223_ ( .A1(_1326_ ), .A2(_1330_ ), .ZN(_1331_ ) );
OAI21_X1 _2224_ ( .A(_1322_ ), .B1(_1331_ ), .B2(_1279_ ), .ZN(_1332_ ) );
AND3_X1 _2225_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(\io_in_a[7] ), .ZN(_1333_ ) );
AND3_X1 _2226_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(\io_in_a[6] ), .ZN(_1334_ ) );
MUX2_X1 _2227_ ( .A(_1333_ ), .B(_1334_ ), .S(_1204_ ), .Z(_1335_ ) );
AND3_X1 _2228_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(\io_in_a[5] ), .ZN(_1336_ ) );
BUF_X4 _2229_ ( .A(_1247_ ), .Z(_1337_ ) );
BUF_X8 _2230_ ( .A(_1337_ ), .Z(_1338_ ) );
BUF_X4 _2231_ ( .A(_1253_ ), .Z(_1339_ ) );
BUF_X8 _2232_ ( .A(_1339_ ), .Z(_1340_ ) );
AND3_X1 _2233_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[4] ), .ZN(_1341_ ) );
MUX2_X1 _2234_ ( .A(_1336_ ), .B(_1341_ ), .S(_1205_ ), .Z(_1342_ ) );
MUX2_X1 _2235_ ( .A(_1335_ ), .B(_1342_ ), .S(_1211_ ), .Z(_1343_ ) );
AND3_X1 _2236_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[3] ), .ZN(_1344_ ) );
AND3_X1 _2237_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[2] ), .ZN(_1345_ ) );
MUX2_X1 _2238_ ( .A(_1344_ ), .B(_1345_ ), .S(_1205_ ), .Z(_1346_ ) );
AND3_X1 _2239_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[1] ), .ZN(_1347_ ) );
AND3_X1 _2240_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[0] ), .ZN(_1348_ ) );
MUX2_X1 _2241_ ( .A(_1347_ ), .B(_1348_ ), .S(_1205_ ), .Z(_1349_ ) );
MUX2_X1 _2242_ ( .A(_1346_ ), .B(_1349_ ), .S(_1211_ ), .Z(_1350_ ) );
BUF_X4 _2243_ ( .A(_1208_ ), .Z(_1351_ ) );
MUX2_X1 _2244_ ( .A(_1343_ ), .B(_1350_ ), .S(_1351_ ), .Z(_1352_ ) );
MUX2_X1 _2245_ ( .A(_1332_ ), .B(_1352_ ), .S(_1215_ ), .Z(_1353_ ) );
MUX2_X1 _2246_ ( .A(_1307_ ), .B(_1353_ ), .S(_1203_ ), .Z(_1354_ ) );
AND2_X1 _2247_ ( .A1(_1237_ ), .A2(_1221_ ), .ZN(_1355_ ) );
INV_X1 _2248_ ( .A(_1355_ ), .ZN(_1356_ ) );
NOR2_X1 _2249_ ( .A1(_0406_ ), .A2(fanout_net_1 ), .ZN(_1357_ ) );
NOR2_X1 _2250_ ( .A1(_1356_ ), .A2(_1357_ ), .ZN(_1358_ ) );
INV_X1 _2251_ ( .A(_1358_ ), .ZN(_1359_ ) );
BUF_X4 _2252_ ( .A(_1308_ ), .Z(_1360_ ) );
BUF_X4 _2253_ ( .A(_1311_ ), .Z(_1361_ ) );
NAND3_X1 _2254_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1022_ ), .ZN(_1362_ ) );
BUF_X4 _2255_ ( .A(_1296_ ), .Z(_1363_ ) );
OAI211_X1 _2256_ ( .A(fanout_net_3 ), .B(_1362_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1364_ ) );
NAND3_X1 _2257_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1324_ ), .ZN(_1365_ ) );
OAI211_X1 _2258_ ( .A(_1206_ ), .B(_1365_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1366_ ) );
AOI21_X1 _2259_ ( .A(_1318_ ), .B1(_1364_ ), .B2(_1366_ ), .ZN(_1367_ ) );
INV_X1 _2260_ ( .A(\io_in_a[13] ), .ZN(_1368_ ) );
NAND3_X2 _2261_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(_1368_ ), .ZN(_1369_ ) );
OAI211_X1 _2262_ ( .A(fanout_net_3 ), .B(_1369_ ), .C1(_1297_ ), .C2(fanout_net_1 ), .ZN(_1370_ ) );
BUF_X16 _2263_ ( .A(_1338_ ), .Z(_1371_ ) );
BUF_X16 _2264_ ( .A(_1340_ ), .Z(_1372_ ) );
NAND3_X2 _2265_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(_1017_ ), .ZN(_1373_ ) );
OAI211_X1 _2266_ ( .A(_1206_ ), .B(_1373_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1374_ ) );
AOI21_X1 _2267_ ( .A(fanout_net_6 ), .B1(_1370_ ), .B2(_1374_ ), .ZN(_1375_ ) );
OAI21_X1 _2268_ ( .A(fanout_net_9 ), .B1(_1367_ ), .B2(_1375_ ), .ZN(_1376_ ) );
NAND3_X1 _2269_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_0994_ ), .ZN(_1377_ ) );
BUF_X4 _2270_ ( .A(_1296_ ), .Z(_1378_ ) );
OAI211_X1 _2271_ ( .A(fanout_net_3 ), .B(_1377_ ), .C1(_1378_ ), .C2(fanout_net_1 ), .ZN(_1379_ ) );
NAND3_X1 _2272_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(_1012_ ), .ZN(_1380_ ) );
OAI211_X1 _2273_ ( .A(_1259_ ), .B(_1380_ ), .C1(_1378_ ), .C2(fanout_net_1 ), .ZN(_1381_ ) );
AOI21_X1 _2274_ ( .A(_1318_ ), .B1(_1379_ ), .B2(_1381_ ), .ZN(_1382_ ) );
INV_X1 _2275_ ( .A(\io_in_a[9] ), .ZN(_1383_ ) );
NAND3_X2 _2276_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(_1383_ ), .ZN(_1384_ ) );
OAI211_X1 _2277_ ( .A(fanout_net_3 ), .B(_1384_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1385_ ) );
BUF_X4 _2278_ ( .A(_1309_ ), .Z(_1386_ ) );
BUF_X4 _2279_ ( .A(_1312_ ), .Z(_1387_ ) );
NAND3_X1 _2280_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_0941_ ), .ZN(_1388_ ) );
OAI211_X1 _2281_ ( .A(_1206_ ), .B(_1388_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1389_ ) );
AOI21_X1 _2282_ ( .A(fanout_net_6 ), .B1(_1385_ ), .B2(_1389_ ), .ZN(_1390_ ) );
OAI21_X1 _2283_ ( .A(_1321_ ), .B1(_1382_ ), .B2(_1390_ ), .ZN(_1391_ ) );
AND2_X1 _2284_ ( .A1(_1376_ ), .A2(_1391_ ), .ZN(_1392_ ) );
NAND3_X1 _2285_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_0332_ ), .ZN(_1393_ ) );
OAI211_X1 _2286_ ( .A(fanout_net_3 ), .B(_1393_ ), .C1(_1378_ ), .C2(fanout_net_1 ), .ZN(_1394_ ) );
NAND3_X1 _2287_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_0471_ ), .ZN(_1395_ ) );
OAI211_X2 _2288_ ( .A(_1259_ ), .B(_1395_ ), .C1(_1378_ ), .C2(fanout_net_1 ), .ZN(_1396_ ) );
AOI21_X1 _2289_ ( .A(_1291_ ), .B1(_1394_ ), .B2(_1396_ ), .ZN(_1397_ ) );
INV_X1 _2290_ ( .A(\io_in_a[5] ), .ZN(_1398_ ) );
NAND3_X1 _2291_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_1398_ ), .ZN(_1399_ ) );
OAI211_X1 _2292_ ( .A(fanout_net_3 ), .B(_1399_ ), .C1(_1378_ ), .C2(fanout_net_1 ), .ZN(_1400_ ) );
NAND3_X1 _2293_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_0385_ ), .ZN(_1401_ ) );
BUF_X4 _2294_ ( .A(_1255_ ), .Z(_1402_ ) );
OAI211_X1 _2295_ ( .A(_1259_ ), .B(_1401_ ), .C1(_1402_ ), .C2(fanout_net_1 ), .ZN(_1403_ ) );
AOI21_X1 _2296_ ( .A(fanout_net_6 ), .B1(_1400_ ), .B2(_1403_ ), .ZN(_1404_ ) );
NOR2_X1 _2297_ ( .A1(_1397_ ), .A2(_1404_ ), .ZN(_1405_ ) );
NAND3_X1 _2298_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_0535_ ), .ZN(_1406_ ) );
OAI211_X1 _2299_ ( .A(fanout_net_3 ), .B(_1406_ ), .C1(_1297_ ), .C2(fanout_net_1 ), .ZN(_1407_ ) );
NAND3_X1 _2300_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(_0503_ ), .ZN(_1408_ ) );
OAI211_X2 _2301_ ( .A(_1206_ ), .B(_1408_ ), .C1(_1297_ ), .C2(fanout_net_1 ), .ZN(_1409_ ) );
AOI21_X1 _2302_ ( .A(_1318_ ), .B1(_1407_ ), .B2(_1409_ ), .ZN(_1410_ ) );
OR4_X1 _2303_ ( .A1(\io_in_b[28] ), .A2(_1244_ ), .A3(_1246_ ), .A4(\io_in_b[25] ), .ZN(_1411_ ) );
OR4_X1 _2304_ ( .A1(\io_in_b[27] ), .A2(_1250_ ), .A3(_1252_ ), .A4(\io_in_b[26] ), .ZN(_1412_ ) );
NOR3_X1 _2305_ ( .A1(_1411_ ), .A2(_1412_ ), .A3(\io_in_a[1] ), .ZN(_1413_ ) );
AOI22_X1 _2306_ ( .A1(_1413_ ), .A2(fanout_net_4 ), .B1(_1256_ ), .B2(_1082_ ), .ZN(_1414_ ) );
NAND3_X1 _2307_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1220_ ), .ZN(_1415_ ) );
AND3_X1 _2308_ ( .A1(_1414_ ), .A2(_1240_ ), .A3(_1415_ ), .ZN(_1416_ ) );
NOR2_X1 _2309_ ( .A1(_1410_ ), .A2(_1416_ ), .ZN(_1417_ ) );
MUX2_X1 _2310_ ( .A(_1405_ ), .B(_1417_ ), .S(_1284_ ), .Z(_1418_ ) );
MUX2_X2 _2311_ ( .A(_1392_ ), .B(_1418_ ), .S(_1283_ ), .Z(_1419_ ) );
NOR2_X1 _2312_ ( .A1(\io_in_b[5] ), .A2(\io_in_b[4] ), .ZN(_1420_ ) );
BUF_X2 _2313_ ( .A(_1420_ ), .Z(_1421_ ) );
AOI21_X1 _2314_ ( .A(_1359_ ), .B1(_1419_ ), .B2(_1421_ ), .ZN(_1422_ ) );
NAND3_X2 _2315_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(_1087_ ), .ZN(_1423_ ) );
OAI211_X1 _2316_ ( .A(fanout_net_4 ), .B(_1423_ ), .C1(_1285_ ), .C2(fanout_net_1 ), .ZN(_1424_ ) );
BUF_X4 _2317_ ( .A(_1204_ ), .Z(_1425_ ) );
NAND3_X1 _2318_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(_1084_ ), .ZN(_1426_ ) );
OAI211_X1 _2319_ ( .A(_1425_ ), .B(_1426_ ), .C1(_1296_ ), .C2(fanout_net_1 ), .ZN(_1427_ ) );
AND2_X1 _2320_ ( .A1(_1424_ ), .A2(_1427_ ), .ZN(_1428_ ) );
OR2_X4 _2321_ ( .A1(_1255_ ), .A2(fanout_net_1 ), .ZN(_1429_ ) );
NAND3_X1 _2322_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(_1091_ ), .ZN(_1430_ ) );
AND2_X1 _2323_ ( .A1(_1429_ ), .A2(_1430_ ), .ZN(_1431_ ) );
AOI21_X1 _2324_ ( .A(_1270_ ), .B1(_1431_ ), .B2(_1259_ ), .ZN(_1432_ ) );
MUX2_X1 _2325_ ( .A(_1428_ ), .B(_1432_ ), .S(fanout_net_6 ), .Z(_1433_ ) );
NAND2_X1 _2326_ ( .A1(_1433_ ), .A2(fanout_net_9 ), .ZN(_1434_ ) );
NAND3_X1 _2327_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(_1063_ ), .ZN(_1435_ ) );
OAI211_X1 _2328_ ( .A(fanout_net_4 ), .B(_1435_ ), .C1(_1285_ ), .C2(fanout_net_1 ), .ZN(_1436_ ) );
NAND3_X1 _2329_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(_1065_ ), .ZN(_1437_ ) );
OAI211_X1 _2330_ ( .A(_1425_ ), .B(_1437_ ), .C1(_1296_ ), .C2(fanout_net_1 ), .ZN(_1438_ ) );
AOI21_X1 _2331_ ( .A(_1291_ ), .B1(_1436_ ), .B2(_1438_ ), .ZN(_1439_ ) );
NAND3_X1 _2332_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(_1069_ ), .ZN(_1440_ ) );
OAI211_X1 _2333_ ( .A(fanout_net_4 ), .B(_1440_ ), .C1(_1402_ ), .C2(fanout_net_1 ), .ZN(_1441_ ) );
NAND3_X4 _2334_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(_1067_ ), .ZN(_1442_ ) );
OAI211_X2 _2335_ ( .A(_1275_ ), .B(_1442_ ), .C1(_1402_ ), .C2(fanout_net_1 ), .ZN(_1443_ ) );
AOI21_X2 _2336_ ( .A(fanout_net_6 ), .B1(_1441_ ), .B2(_1443_ ), .ZN(_1444_ ) );
OR3_X4 _2337_ ( .A1(_1439_ ), .A2(_1444_ ), .A3(fanout_net_9 ), .ZN(_1445_ ) );
NAND3_X1 _2338_ ( .A1(_1434_ ), .A2(fanout_net_12 ), .A3(_1445_ ), .ZN(_1446_ ) );
NAND3_X2 _2339_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(_1048_ ), .ZN(_1447_ ) );
OAI211_X1 _2340_ ( .A(fanout_net_4 ), .B(_1447_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1448_ ) );
NAND3_X1 _2341_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1033_ ), .ZN(_1449_ ) );
OAI211_X1 _2342_ ( .A(_1259_ ), .B(_1449_ ), .C1(_1378_ ), .C2(fanout_net_1 ), .ZN(_1450_ ) );
AOI21_X1 _2343_ ( .A(_1212_ ), .B1(_1448_ ), .B2(_1450_ ), .ZN(_1451_ ) );
INV_X1 _2344_ ( .A(\io_in_a[21] ), .ZN(_1452_ ) );
NAND3_X1 _2345_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1452_ ), .ZN(_1453_ ) );
OAI211_X1 _2346_ ( .A(fanout_net_4 ), .B(_1453_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1454_ ) );
NAND3_X2 _2347_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(_1028_ ), .ZN(_1455_ ) );
OAI211_X1 _2348_ ( .A(_1206_ ), .B(_1455_ ), .C1(_1363_ ), .C2(fanout_net_1 ), .ZN(_1456_ ) );
AOI21_X1 _2349_ ( .A(fanout_net_6 ), .B1(_1454_ ), .B2(_1456_ ), .ZN(_1457_ ) );
OAI21_X1 _2350_ ( .A(fanout_net_9 ), .B1(_1451_ ), .B2(_1457_ ), .ZN(_1458_ ) );
NAND3_X1 _2351_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1041_ ), .ZN(_1459_ ) );
OAI211_X1 _2352_ ( .A(fanout_net_4 ), .B(_1459_ ), .C1(_1378_ ), .C2(fanout_net_2 ), .ZN(_1460_ ) );
NAND3_X1 _2353_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1043_ ), .ZN(_1461_ ) );
OAI211_X1 _2354_ ( .A(_1259_ ), .B(_1461_ ), .C1(_1378_ ), .C2(fanout_net_2 ), .ZN(_1462_ ) );
AOI21_X1 _2355_ ( .A(_1212_ ), .B1(_1460_ ), .B2(_1462_ ), .ZN(_1463_ ) );
INV_X1 _2356_ ( .A(\io_in_a[17] ), .ZN(_1464_ ) );
NAND3_X1 _2357_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1464_ ), .ZN(_1465_ ) );
OAI211_X1 _2358_ ( .A(fanout_net_4 ), .B(_1465_ ), .C1(_1297_ ), .C2(fanout_net_2 ), .ZN(_1466_ ) );
NAND3_X1 _2359_ ( .A1(_1360_ ), .A2(_1361_ ), .A3(_1035_ ), .ZN(_1467_ ) );
OAI211_X1 _2360_ ( .A(_1206_ ), .B(_1467_ ), .C1(_1297_ ), .C2(fanout_net_2 ), .ZN(_1468_ ) );
AOI21_X1 _2361_ ( .A(fanout_net_6 ), .B1(_1466_ ), .B2(_1468_ ), .ZN(_1469_ ) );
OAI21_X1 _2362_ ( .A(_1284_ ), .B1(_1463_ ), .B2(_1469_ ), .ZN(_1470_ ) );
AND2_X1 _2363_ ( .A1(_1458_ ), .A2(_1470_ ), .ZN(_1471_ ) );
OR2_X1 _2364_ ( .A1(_1471_ ), .A2(fanout_net_12 ), .ZN(_1472_ ) );
NOR2_X1 _2365_ ( .A1(_1202_ ), .A2(\io_in_b[5] ), .ZN(_1473_ ) );
BUF_X2 _2366_ ( .A(_1473_ ), .Z(_1474_ ) );
NAND3_X1 _2367_ ( .A1(_1446_ ), .A2(_1472_ ), .A3(_1474_ ), .ZN(_1475_ ) );
AOI22_X1 _2368_ ( .A1(_1239_ ), .A2(_1354_ ), .B1(_1422_ ), .B2(_1475_ ), .ZN(_1476_ ) );
AOI21_X2 _2369_ ( .A(_1088_ ), .B1(_1073_ ), .B2(_1080_ ), .ZN(_1477_ ) );
NOR2_X1 _2370_ ( .A1(_1477_ ), .A2(_1074_ ), .ZN(_1478_ ) );
NOR2_X1 _2371_ ( .A1(_1091_ ), .A2(\io_in_b[30] ), .ZN(_1479_ ) );
NOR2_X2 _2372_ ( .A1(_1478_ ), .A2(_1479_ ), .ZN(_1480_ ) );
INV_X1 _2373_ ( .A(_1480_ ), .ZN(_1481_ ) );
NOR2_X4 _2374_ ( .A1(_1090_ ), .A2(_1092_ ), .ZN(_1482_ ) );
MUX2_X2 _2375_ ( .A(_1481_ ), .B(_1482_ ), .S(_0052_ ), .Z(_1483_ ) );
BUF_X4 _2376_ ( .A(_1226_ ), .Z(_1484_ ) );
NAND3_X1 _2377_ ( .A1(_1484_ ), .A2(\io_sw[3] ), .A3(_1094_ ), .ZN(_1485_ ) );
OAI211_X1 _2378_ ( .A(_1236_ ), .B(_1476_ ), .C1(_1483_ ), .C2(_1485_ ), .ZN(\io_out[0] ) );
XNOR2_X1 _2379_ ( .A(_1480_ ), .B(_0062_ ), .ZN(_1486_ ) );
BUF_X2 _2380_ ( .A(_1098_ ), .Z(_1487_ ) );
NAND2_X1 _2381_ ( .A1(_1486_ ), .A2(_1487_ ), .ZN(_1488_ ) );
NAND2_X4 _2382_ ( .A1(_1189_ ), .A2(_1193_ ), .ZN(_1489_ ) );
NAND2_X4 _2383_ ( .A1(_1489_ ), .A2(_1074_ ), .ZN(_1490_ ) );
NAND2_X2 _2384_ ( .A1(_1490_ ), .A2(_1196_ ), .ZN(_1491_ ) );
XNOR2_X1 _2385_ ( .A(_1491_ ), .B(_0062_ ), .ZN(_1492_ ) );
NAND2_X1 _2386_ ( .A1(_1492_ ), .A2(_1106_ ), .ZN(_1493_ ) );
NOR2_X1 _2387_ ( .A1(_1082_ ), .A2(fanout_net_4 ), .ZN(_1494_ ) );
AND3_X1 _2388_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1494_ ), .ZN(_1495_ ) );
BUF_X4 _2389_ ( .A(_1351_ ), .Z(_1496_ ) );
BUF_X2 _2390_ ( .A(_1496_ ), .Z(_1497_ ) );
BUF_X2 _2391_ ( .A(_1327_ ), .Z(_1498_ ) );
AND3_X1 _2392_ ( .A1(_1495_ ), .A2(_1497_ ), .A3(_1498_ ), .ZN(_1499_ ) );
BUF_X4 _2393_ ( .A(_1215_ ), .Z(_1500_ ) );
BUF_X2 _2394_ ( .A(_1500_ ), .Z(_1501_ ) );
AND2_X1 _2395_ ( .A1(_1238_ ), .A2(_1420_ ), .ZN(_1502_ ) );
BUF_X2 _2396_ ( .A(_1502_ ), .Z(_1503_ ) );
NAND3_X1 _2397_ ( .A1(_1499_ ), .A2(_1501_ ), .A3(_1503_ ), .ZN(_1504_ ) );
AND2_X2 _2398_ ( .A1(_1218_ ), .A2(_1202_ ), .ZN(_1505_ ) );
BUF_X2 _2399_ ( .A(_1505_ ), .Z(_1506_ ) );
BUF_X2 _2400_ ( .A(_1506_ ), .Z(_1507_ ) );
AND2_X1 _2401_ ( .A1(fanout_net_4 ), .A2(\io_in_a[26] ), .ZN(_1508_ ) );
INV_X1 _2402_ ( .A(_1508_ ), .ZN(_1509_ ) );
BUF_X4 _2403_ ( .A(_1327_ ), .Z(_1510_ ) );
OAI211_X1 _2404_ ( .A(_1509_ ), .B(_1510_ ), .C1(fanout_net_4 ), .C2(_1063_ ), .ZN(_1511_ ) );
NOR2_X1 _2405_ ( .A1(_1069_ ), .A2(fanout_net_4 ), .ZN(_1512_ ) );
INV_X1 _2406_ ( .A(_1512_ ), .ZN(_1513_ ) );
AND2_X1 _2407_ ( .A1(fanout_net_4 ), .A2(\io_in_a[24] ), .ZN(_1514_ ) );
INV_X1 _2408_ ( .A(_1514_ ), .ZN(_1515_ ) );
NAND3_X1 _2409_ ( .A1(_1513_ ), .A2(fanout_net_6 ), .A3(_1515_ ), .ZN(_1516_ ) );
NAND3_X1 _2410_ ( .A1(_1511_ ), .A2(_1516_ ), .A3(fanout_net_9 ), .ZN(_1517_ ) );
BUF_X4 _2411_ ( .A(_1284_ ), .Z(_1518_ ) );
NAND2_X1 _2412_ ( .A1(fanout_net_4 ), .A2(\io_in_a[30] ), .ZN(_1519_ ) );
OAI211_X1 _2413_ ( .A(_1519_ ), .B(_1498_ ), .C1(fanout_net_4 ), .C2(_1082_ ), .ZN(_1520_ ) );
NAND2_X1 _2414_ ( .A1(_1204_ ), .A2(\io_in_a[29] ), .ZN(_1521_ ) );
NAND2_X1 _2415_ ( .A1(fanout_net_4 ), .A2(\io_in_a[28] ), .ZN(_1522_ ) );
NAND2_X1 _2416_ ( .A1(_1521_ ), .A2(_1522_ ), .ZN(_1523_ ) );
OAI211_X1 _2417_ ( .A(_1518_ ), .B(_1520_ ), .C1(_1523_ ), .C2(_1498_ ), .ZN(_1524_ ) );
AOI21_X1 _2418_ ( .A(fanout_net_12 ), .B1(_1517_ ), .B2(_1524_ ), .ZN(_1525_ ) );
NOR2_X1 _2419_ ( .A1(_1452_ ), .A2(fanout_net_4 ), .ZN(_1526_ ) );
AND2_X1 _2420_ ( .A1(fanout_net_4 ), .A2(\io_in_a[20] ), .ZN(_1527_ ) );
OR3_X1 _2421_ ( .A1(_1526_ ), .A2(_1527_ ), .A3(_1327_ ), .ZN(_1528_ ) );
NOR2_X1 _2422_ ( .A1(_1048_ ), .A2(fanout_net_4 ), .ZN(_1529_ ) );
INV_X1 _2423_ ( .A(_1529_ ), .ZN(_1530_ ) );
AND2_X1 _2424_ ( .A1(fanout_net_4 ), .A2(\io_in_a[22] ), .ZN(_1531_ ) );
INV_X1 _2425_ ( .A(_1531_ ), .ZN(_1532_ ) );
NAND3_X1 _2426_ ( .A1(_1530_ ), .A2(_1510_ ), .A3(_1532_ ), .ZN(_1533_ ) );
NAND2_X1 _2427_ ( .A1(_1528_ ), .A2(_1533_ ), .ZN(_1534_ ) );
BUF_X4 _2428_ ( .A(_1321_ ), .Z(_1535_ ) );
NAND2_X1 _2429_ ( .A1(_1534_ ), .A2(_1535_ ), .ZN(_1536_ ) );
NOR2_X1 _2430_ ( .A1(_1041_ ), .A2(fanout_net_4 ), .ZN(_1537_ ) );
AND2_X1 _2431_ ( .A1(fanout_net_4 ), .A2(\io_in_a[18] ), .ZN(_1538_ ) );
OAI21_X1 _2432_ ( .A(_0589_ ), .B1(_1537_ ), .B2(_1538_ ), .ZN(_1539_ ) );
NOR2_X1 _2433_ ( .A1(_1464_ ), .A2(fanout_net_4 ), .ZN(_1540_ ) );
AND2_X1 _2434_ ( .A1(fanout_net_4 ), .A2(\io_in_a[16] ), .ZN(_1541_ ) );
OAI21_X1 _2435_ ( .A(fanout_net_6 ), .B1(_1540_ ), .B2(_1541_ ), .ZN(_1542_ ) );
NAND3_X1 _2436_ ( .A1(_1539_ ), .A2(_1542_ ), .A3(fanout_net_9 ), .ZN(_1543_ ) );
AND3_X1 _2437_ ( .A1(_1536_ ), .A2(fanout_net_12 ), .A3(_1543_ ), .ZN(_1544_ ) );
OAI21_X1 _2438_ ( .A(_1507_ ), .B1(_1525_ ), .B2(_1544_ ), .ZN(_1545_ ) );
NOR2_X1 _2439_ ( .A1(_0994_ ), .A2(fanout_net_4 ), .ZN(_1546_ ) );
AND2_X1 _2440_ ( .A1(fanout_net_4 ), .A2(\io_in_a[10] ), .ZN(_1547_ ) );
OAI21_X1 _2441_ ( .A(_1290_ ), .B1(_1546_ ), .B2(_1547_ ), .ZN(_1548_ ) );
NOR2_X1 _2442_ ( .A1(_1383_ ), .A2(fanout_net_4 ), .ZN(_1549_ ) );
AND2_X1 _2443_ ( .A1(fanout_net_4 ), .A2(\io_in_a[8] ), .ZN(_1550_ ) );
OAI21_X1 _2444_ ( .A(fanout_net_6 ), .B1(_1549_ ), .B2(_1550_ ), .ZN(_1551_ ) );
NAND2_X1 _2445_ ( .A1(_1548_ ), .A2(_1551_ ), .ZN(_1552_ ) );
NAND2_X1 _2446_ ( .A1(_1552_ ), .A2(fanout_net_9 ), .ZN(_1553_ ) );
NOR2_X1 _2447_ ( .A1(_1022_ ), .A2(fanout_net_4 ), .ZN(_1554_ ) );
AND2_X1 _2448_ ( .A1(fanout_net_4 ), .A2(\io_in_a[14] ), .ZN(_1555_ ) );
OR3_X1 _2449_ ( .A1(_1554_ ), .A2(_1555_ ), .A3(fanout_net_6 ), .ZN(_1556_ ) );
NOR2_X1 _2450_ ( .A1(_1368_ ), .A2(fanout_net_5 ), .ZN(_1557_ ) );
INV_X1 _2451_ ( .A(_1557_ ), .ZN(_1558_ ) );
AND2_X1 _2452_ ( .A1(fanout_net_5 ), .A2(\io_in_a[12] ), .ZN(_1559_ ) );
INV_X1 _2453_ ( .A(_1559_ ), .ZN(_1560_ ) );
NAND3_X1 _2454_ ( .A1(_1558_ ), .A2(fanout_net_6 ), .A3(_1560_ ), .ZN(_1561_ ) );
NAND3_X1 _2455_ ( .A1(_1556_ ), .A2(_1561_ ), .A3(_1535_ ), .ZN(_1562_ ) );
NAND3_X1 _2456_ ( .A1(_1553_ ), .A2(_1562_ ), .A3(_1500_ ), .ZN(_1563_ ) );
AND2_X1 _2457_ ( .A1(_1218_ ), .A2(\io_in_b[4] ), .ZN(_1564_ ) );
BUF_X2 _2458_ ( .A(_1564_ ), .Z(_1565_ ) );
NOR2_X1 _2459_ ( .A1(_0332_ ), .A2(fanout_net_5 ), .ZN(_1566_ ) );
AND2_X1 _2460_ ( .A1(fanout_net_5 ), .A2(\io_in_a[6] ), .ZN(_1567_ ) );
OAI21_X1 _2461_ ( .A(_1210_ ), .B1(_1566_ ), .B2(_1567_ ), .ZN(_1568_ ) );
NOR2_X1 _2462_ ( .A1(_1398_ ), .A2(fanout_net_5 ), .ZN(_1569_ ) );
AND2_X1 _2463_ ( .A1(fanout_net_5 ), .A2(\io_in_a[4] ), .ZN(_1570_ ) );
OAI21_X1 _2464_ ( .A(fanout_net_6 ), .B1(_1569_ ), .B2(_1570_ ), .ZN(_1571_ ) );
AND3_X1 _2465_ ( .A1(_1568_ ), .A2(_1571_ ), .A3(_1208_ ), .ZN(_1572_ ) );
NOR2_X1 _2466_ ( .A1(_0535_ ), .A2(fanout_net_5 ), .ZN(_1573_ ) );
AND2_X1 _2467_ ( .A1(fanout_net_5 ), .A2(\io_in_a[2] ), .ZN(_1574_ ) );
NOR2_X1 _2468_ ( .A1(_1573_ ), .A2(_1574_ ), .ZN(_1575_ ) );
AOI21_X1 _2469_ ( .A(_1123_ ), .B1(_1204_ ), .B2(\io_in_a[1] ), .ZN(_1576_ ) );
MUX2_X1 _2470_ ( .A(_1575_ ), .B(_1576_ ), .S(fanout_net_6 ), .Z(_1577_ ) );
AOI21_X1 _2471_ ( .A(_1572_ ), .B1(_1577_ ), .B2(fanout_net_9 ), .ZN(_1578_ ) );
BUF_X2 _2472_ ( .A(_1283_ ), .Z(_1579_ ) );
OAI211_X1 _2473_ ( .A(_1563_ ), .B(_1565_ ), .C1(_1578_ ), .C2(_1579_ ), .ZN(_1580_ ) );
BUF_X4 _2474_ ( .A(_1223_ ), .Z(_1581_ ) );
BUF_X4 _2475_ ( .A(_1581_ ), .Z(_1582_ ) );
AOI22_X1 _2476_ ( .A1(_0030_ ), .A2(_1228_ ), .B1(_1582_ ), .B2(_0052_ ), .ZN(_1583_ ) );
BUF_X4 _2477_ ( .A(_1232_ ), .Z(_1584_ ) );
BUF_X4 _2478_ ( .A(_1584_ ), .Z(_1585_ ) );
INV_X1 _2479_ ( .A(_0041_ ), .ZN(_1586_ ) );
AOI22_X1 _2480_ ( .A1(_1355_ ), .A2(fanout_net_2 ), .B1(_1585_ ), .B2(_1586_ ), .ZN(_1587_ ) );
AND4_X1 _2481_ ( .A1(_1545_ ), .A2(_1580_ ), .A3(_1583_ ), .A4(_1587_ ), .ZN(_1588_ ) );
NAND4_X1 _2482_ ( .A1(_1488_ ), .A2(_1493_ ), .A3(_1504_ ), .A4(_1588_ ), .ZN(\io_out[31] ) );
AND2_X4 _2483_ ( .A1(_0931_ ), .A2(_1026_ ), .ZN(_1589_ ) );
NOR2_X4 _2484_ ( .A1(_1589_ ), .A2(_0278_ ), .ZN(_1590_ ) );
AND3_X4 _2485_ ( .A1(_1590_ ), .A2(_0245_ ), .A3(_0202_ ), .ZN(_1591_ ) );
NOR2_X4 _2486_ ( .A1(_1591_ ), .A2(_1046_ ), .ZN(_1592_ ) );
NOR2_X4 _2487_ ( .A1(_1592_ ), .A2(_0073_ ), .ZN(_1593_ ) );
NOR2_X1 _2488_ ( .A1(_1028_ ), .A2(\io_in_b[20] ), .ZN(_1594_ ) );
NOR2_X4 _2489_ ( .A1(_1593_ ), .A2(_1594_ ), .ZN(_1595_ ) );
NOR2_X2 _2490_ ( .A1(_1595_ ), .A2(_0084_ ), .ZN(_1596_ ) );
AOI21_X2 _2491_ ( .A(_1596_ ), .B1(\io_in_a[21] ), .B2(_1030_ ), .ZN(_1597_ ) );
NOR2_X2 _2492_ ( .A1(_1597_ ), .A2(_0127_ ), .ZN(_1598_ ) );
INV_X4 _2493_ ( .A(_1598_ ), .ZN(_1599_ ) );
AOI21_X1 _2494_ ( .A(_1101_ ), .B1(_1597_ ), .B2(_0127_ ), .ZN(_1600_ ) );
NOR2_X1 _2495_ ( .A1(_1209_ ), .A2(fanout_net_2 ), .ZN(_1601_ ) );
INV_X1 _2496_ ( .A(_1601_ ), .ZN(_1602_ ) );
NAND2_X1 _2497_ ( .A1(_1432_ ), .A2(_1327_ ), .ZN(_1603_ ) );
NAND2_X1 _2498_ ( .A1(_1082_ ), .A2(fanout_net_6 ), .ZN(_1604_ ) );
AND2_X1 _2499_ ( .A1(_1603_ ), .A2(_1604_ ), .ZN(_1605_ ) );
OAI211_X1 _2500_ ( .A(fanout_net_12 ), .B(_1602_ ), .C1(_1605_ ), .C2(fanout_net_9 ), .ZN(_1606_ ) );
BUF_X2 _2501_ ( .A(_1421_ ), .Z(_1607_ ) );
AOI21_X1 _2502_ ( .A(_1291_ ), .B1(_1441_ ), .B2(_1443_ ), .ZN(_1608_ ) );
AOI21_X1 _2503_ ( .A(fanout_net_6 ), .B1(_1448_ ), .B2(_1450_ ), .ZN(_1609_ ) );
OAI21_X1 _2504_ ( .A(_1518_ ), .B1(_1608_ ), .B2(_1609_ ), .ZN(_1610_ ) );
BUF_X4 _2505_ ( .A(_1210_ ), .Z(_1611_ ) );
NAND3_X1 _2506_ ( .A1(_1436_ ), .A2(_1438_ ), .A3(_1611_ ), .ZN(_1612_ ) );
NAND3_X1 _2507_ ( .A1(_1424_ ), .A2(_1427_ ), .A3(fanout_net_6 ), .ZN(_1613_ ) );
NAND3_X1 _2508_ ( .A1(_1612_ ), .A2(_1613_ ), .A3(fanout_net_9 ), .ZN(_1614_ ) );
NAND2_X1 _2509_ ( .A1(_1610_ ), .A2(_1614_ ), .ZN(_1615_ ) );
NAND2_X1 _2510_ ( .A1(_1615_ ), .A2(_1579_ ), .ZN(_1616_ ) );
NAND3_X1 _2511_ ( .A1(_1606_ ), .A2(_1607_ ), .A3(_1616_ ), .ZN(_1617_ ) );
AOI21_X1 _2512_ ( .A(fanout_net_2 ), .B1(_0406_ ), .B2(_1202_ ), .ZN(_1618_ ) );
NOR2_X1 _2513_ ( .A1(_1356_ ), .A2(_1618_ ), .ZN(_1619_ ) );
AOI22_X1 _2514_ ( .A1(_1599_ ), .A2(_1600_ ), .B1(_1617_ ), .B2(_1619_ ), .ZN(_1620_ ) );
NOR4_X1 _2515_ ( .A1(_1161_ ), .A2(_0245_ ), .A3(_0289_ ), .A4(_1171_ ), .ZN(_1621_ ) );
OAI21_X1 _2516_ ( .A(_1163_ ), .B1(_1621_ ), .B2(_1173_ ), .ZN(_1622_ ) );
AND3_X1 _2517_ ( .A1(_1622_ ), .A2(_0138_ ), .A3(_1177_ ), .ZN(_1623_ ) );
AOI21_X1 _2518_ ( .A(_0138_ ), .B1(_1622_ ), .B2(_1177_ ), .ZN(_1624_ ) );
INV_X1 _2519_ ( .A(_1105_ ), .ZN(_1625_ ) );
BUF_X2 _2520_ ( .A(_1625_ ), .Z(_1626_ ) );
OR3_X1 _2521_ ( .A1(_1623_ ), .A2(_1624_ ), .A3(_1626_ ), .ZN(_1627_ ) );
AOI211_X1 _2522_ ( .A(_1498_ ), .B(_1257_ ), .C1(_1274_ ), .C2(_1276_ ), .ZN(_1628_ ) );
AOI211_X1 _2523_ ( .A(fanout_net_6 ), .B(_1257_ ), .C1(_1258_ ), .C2(_1260_ ), .ZN(_1629_ ) );
OAI21_X1 _2524_ ( .A(fanout_net_9 ), .B1(_1628_ ), .B2(_1629_ ), .ZN(_1630_ ) );
AOI211_X1 _2525_ ( .A(_1498_ ), .B(_1257_ ), .C1(_1263_ ), .C2(_1265_ ), .ZN(_1631_ ) );
OAI21_X1 _2526_ ( .A(_1298_ ), .B1(_1287_ ), .B2(_1288_ ), .ZN(_1632_ ) );
NOR2_X1 _2527_ ( .A1(_1632_ ), .A2(fanout_net_6 ), .ZN(_1633_ ) );
OAI21_X1 _2528_ ( .A(_1518_ ), .B1(_1631_ ), .B2(_1633_ ), .ZN(_1634_ ) );
AOI21_X1 _2529_ ( .A(fanout_net_12 ), .B1(_1630_ ), .B2(_1634_ ), .ZN(_1635_ ) );
BUF_X2 _2530_ ( .A(_1282_ ), .Z(_1636_ ) );
NOR4_X1 _2531_ ( .A1(_1272_ ), .A2(_1636_ ), .A3(fanout_net_9 ), .A4(fanout_net_6 ), .ZN(_1637_ ) );
OAI21_X1 _2532_ ( .A(_1503_ ), .B1(_1635_ ), .B2(_1637_ ), .ZN(_1638_ ) );
OAI21_X1 _2533_ ( .A(_1510_ ), .B1(_1287_ ), .B2(_1292_ ), .ZN(_1639_ ) );
OAI21_X1 _2534_ ( .A(fanout_net_6 ), .B1(_1293_ ), .B2(_1299_ ), .ZN(_1640_ ) );
NAND2_X1 _2535_ ( .A1(_1639_ ), .A2(_1640_ ), .ZN(_1641_ ) );
NAND2_X1 _2536_ ( .A1(_1641_ ), .A2(_1535_ ), .ZN(_1642_ ) );
OAI21_X1 _2537_ ( .A(_1510_ ), .B1(_1300_ ), .B2(_1302_ ), .ZN(_1643_ ) );
OAI21_X1 _2538_ ( .A(fanout_net_6 ), .B1(_1303_ ), .B2(_1323_ ), .ZN(_1644_ ) );
NAND2_X1 _2539_ ( .A1(_1643_ ), .A2(_1644_ ), .ZN(_1645_ ) );
NAND2_X1 _2540_ ( .A1(_1645_ ), .A2(fanout_net_9 ), .ZN(_1646_ ) );
BUF_X4 _2541_ ( .A(_1283_ ), .Z(_1647_ ) );
NAND3_X1 _2542_ ( .A1(_1642_ ), .A2(_1646_ ), .A3(_1647_ ), .ZN(_1648_ ) );
OAI21_X1 _2543_ ( .A(_1611_ ), .B1(_1325_ ), .B2(_1328_ ), .ZN(_1649_ ) );
AND2_X1 _2544_ ( .A1(fanout_net_5 ), .A2(\io_in_a[11] ), .ZN(_1650_ ) );
OAI21_X1 _2545_ ( .A(fanout_net_6 ), .B1(_1329_ ), .B2(_1650_ ), .ZN(_1651_ ) );
NAND2_X1 _2546_ ( .A1(_1649_ ), .A2(_1651_ ), .ZN(_1652_ ) );
NAND2_X1 _2547_ ( .A1(_1652_ ), .A2(_1351_ ), .ZN(_1653_ ) );
NOR2_X1 _2548_ ( .A1(_0941_ ), .A2(fanout_net_5 ), .ZN(_1654_ ) );
AND2_X1 _2549_ ( .A1(fanout_net_5 ), .A2(\io_in_a[7] ), .ZN(_1655_ ) );
OR3_X1 _2550_ ( .A1(_1654_ ), .A2(_1655_ ), .A3(_1290_ ), .ZN(_1656_ ) );
NOR2_X1 _2551_ ( .A1(_1012_ ), .A2(fanout_net_5 ), .ZN(_1657_ ) );
AND2_X1 _2552_ ( .A1(fanout_net_5 ), .A2(\io_in_a[9] ), .ZN(_1658_ ) );
OR3_X1 _2553_ ( .A1(_1657_ ), .A2(_1658_ ), .A3(fanout_net_7 ), .ZN(_1659_ ) );
NAND3_X1 _2554_ ( .A1(_1656_ ), .A2(_1659_ ), .A3(fanout_net_9 ), .ZN(_1660_ ) );
NAND3_X1 _2555_ ( .A1(_1653_ ), .A2(_1660_ ), .A3(fanout_net_12 ), .ZN(_1661_ ) );
NAND3_X1 _2556_ ( .A1(_1648_ ), .A2(_1661_ ), .A3(_1507_ ), .ZN(_1662_ ) );
NOR2_X1 _2557_ ( .A1(_0503_ ), .A2(fanout_net_5 ), .ZN(_1663_ ) );
AND2_X1 _2558_ ( .A1(fanout_net_5 ), .A2(\io_in_a[1] ), .ZN(_1664_ ) );
OAI21_X1 _2559_ ( .A(_1210_ ), .B1(_1663_ ), .B2(_1664_ ), .ZN(_1665_ ) );
NAND3_X1 _2560_ ( .A1(_1425_ ), .A2(\io_in_a[0] ), .A3(fanout_net_7 ), .ZN(_1666_ ) );
NAND2_X1 _2561_ ( .A1(_1665_ ), .A2(_1666_ ), .ZN(_1667_ ) );
NOR2_X1 _2562_ ( .A1(_0471_ ), .A2(fanout_net_5 ), .ZN(_1668_ ) );
AND2_X1 _2563_ ( .A1(fanout_net_5 ), .A2(\io_in_a[5] ), .ZN(_1669_ ) );
OAI21_X1 _2564_ ( .A(_1210_ ), .B1(_1668_ ), .B2(_1669_ ), .ZN(_1670_ ) );
NOR2_X1 _2565_ ( .A1(_0385_ ), .A2(fanout_net_5 ), .ZN(_1671_ ) );
AND2_X1 _2566_ ( .A1(fanout_net_5 ), .A2(\io_in_a[3] ), .ZN(_1672_ ) );
OAI21_X1 _2567_ ( .A(fanout_net_7 ), .B1(_1671_ ), .B2(_1672_ ), .ZN(_1673_ ) );
NAND2_X1 _2568_ ( .A1(_1670_ ), .A2(_1673_ ), .ZN(_1674_ ) );
MUX2_X1 _2569_ ( .A(_1667_ ), .B(_1674_ ), .S(_1208_ ), .Z(_1675_ ) );
BUF_X4 _2570_ ( .A(_1215_ ), .Z(_1676_ ) );
BUF_X4 _2571_ ( .A(_1676_ ), .Z(_1677_ ) );
NAND3_X1 _2572_ ( .A1(_1675_ ), .A2(_1677_ ), .A3(_1565_ ), .ZN(_1678_ ) );
OAI21_X1 _2573_ ( .A(_1585_ ), .B1(\io_in_a[22] ), .B2(\io_in_b[22] ), .ZN(_1679_ ) );
AOI22_X1 _2574_ ( .A1(_1180_ ), .A2(_1228_ ), .B1(_1582_ ), .B2(_0127_ ), .ZN(_1680_ ) );
AND4_X1 _2575_ ( .A1(_1662_ ), .A2(_1678_ ), .A3(_1679_ ), .A4(_1680_ ), .ZN(_1681_ ) );
NAND4_X1 _2576_ ( .A1(_1620_ ), .A2(_1627_ ), .A3(_1638_ ), .A4(_1681_ ), .ZN(\io_out[22] ) );
AND2_X1 _2577_ ( .A1(_1595_ ), .A2(_0084_ ), .ZN(_1682_ ) );
OR3_X1 _2578_ ( .A1(_1682_ ), .A2(_1596_ ), .A3(_1100_ ), .ZN(_1683_ ) );
OR2_X1 _2579_ ( .A1(_1621_ ), .A2(_1173_ ), .ZN(_1684_ ) );
AOI21_X1 _2580_ ( .A(_1176_ ), .B1(_1684_ ), .B2(_0073_ ), .ZN(_1685_ ) );
XNOR2_X1 _2581_ ( .A(_1685_ ), .B(_0084_ ), .ZN(_1686_ ) );
AND2_X1 _2582_ ( .A1(_1686_ ), .A2(_1106_ ), .ZN(_1687_ ) );
INV_X1 _2583_ ( .A(_1502_ ), .ZN(_1688_ ) );
AOI211_X1 _2584_ ( .A(fanout_net_7 ), .B(_1257_ ), .C1(_1519_ ), .C2(_1521_ ), .ZN(_1689_ ) );
AND4_X1 _2585_ ( .A1(fanout_net_7 ), .A2(_1309_ ), .A3(_1312_ ), .A4(_1494_ ), .ZN(_1690_ ) );
OAI211_X1 _2586_ ( .A(fanout_net_12 ), .B(_1497_ ), .C1(_1689_ ), .C2(_1690_ ), .ZN(_1691_ ) );
OAI211_X1 _2587_ ( .A(_1285_ ), .B(fanout_net_7 ), .C1(_1514_ ), .C2(_1529_ ), .ZN(_1692_ ) );
OAI211_X1 _2588_ ( .A(_1285_ ), .B(_1210_ ), .C1(_1526_ ), .C2(_1531_ ), .ZN(_1693_ ) );
AOI21_X1 _2589_ ( .A(fanout_net_9 ), .B1(_1692_ ), .B2(_1693_ ), .ZN(_1694_ ) );
OAI211_X1 _2590_ ( .A(_1285_ ), .B(_1210_ ), .C1(_1512_ ), .C2(_1508_ ), .ZN(_1695_ ) );
OAI21_X1 _2591_ ( .A(_1522_ ), .B1(_1063_ ), .B2(fanout_net_5 ), .ZN(_1696_ ) );
NAND4_X1 _2592_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(fanout_net_7 ), .A4(_1696_ ), .ZN(_1697_ ) );
AOI21_X1 _2593_ ( .A(_1279_ ), .B1(_1695_ ), .B2(_1697_ ), .ZN(_1698_ ) );
OAI21_X1 _2594_ ( .A(_1216_ ), .B1(_1694_ ), .B2(_1698_ ), .ZN(_1699_ ) );
AOI21_X1 _2595_ ( .A(_1688_ ), .B1(_1691_ ), .B2(_1699_ ), .ZN(_1700_ ) );
OR3_X1 _2596_ ( .A1(_1566_ ), .A2(_1567_ ), .A3(_1290_ ), .ZN(_1701_ ) );
OR3_X1 _2597_ ( .A1(_1549_ ), .A2(_1550_ ), .A3(fanout_net_7 ), .ZN(_1702_ ) );
NAND3_X1 _2598_ ( .A1(_1701_ ), .A2(_1702_ ), .A3(fanout_net_9 ), .ZN(_1703_ ) );
OR3_X1 _2599_ ( .A1(_1546_ ), .A2(_1547_ ), .A3(_1210_ ), .ZN(_1704_ ) );
NAND3_X1 _2600_ ( .A1(_1558_ ), .A2(_1211_ ), .A3(_1560_ ), .ZN(_1705_ ) );
NAND3_X1 _2601_ ( .A1(_1704_ ), .A2(_1705_ ), .A3(_1496_ ), .ZN(_1706_ ) );
AOI21_X1 _2602_ ( .A(_1636_ ), .B1(_1703_ ), .B2(_1706_ ), .ZN(_1707_ ) );
OAI21_X1 _2603_ ( .A(_1327_ ), .B1(_1526_ ), .B2(_1527_ ), .ZN(_1708_ ) );
OAI21_X1 _2604_ ( .A(fanout_net_7 ), .B1(_1537_ ), .B2(_1538_ ), .ZN(_1709_ ) );
AOI21_X1 _2605_ ( .A(fanout_net_9 ), .B1(_1708_ ), .B2(_1709_ ), .ZN(_1710_ ) );
OAI21_X1 _2606_ ( .A(_1290_ ), .B1(_1540_ ), .B2(_1541_ ), .ZN(_1711_ ) );
OAI21_X1 _2607_ ( .A(fanout_net_7 ), .B1(_1554_ ), .B2(_1555_ ), .ZN(_1712_ ) );
AOI21_X1 _2608_ ( .A(_1284_ ), .B1(_1711_ ), .B2(_1712_ ), .ZN(_1713_ ) );
OR2_X1 _2609_ ( .A1(_1710_ ), .A2(_1713_ ), .ZN(_1714_ ) );
AOI21_X1 _2610_ ( .A(_1707_ ), .B1(_1216_ ), .B2(_1714_ ), .ZN(_1715_ ) );
INV_X1 _2611_ ( .A(_1505_ ), .ZN(_1716_ ) );
NOR2_X1 _2612_ ( .A1(_1715_ ), .A2(_1716_ ), .ZN(_1717_ ) );
OAI21_X1 _2613_ ( .A(_1211_ ), .B1(_1569_ ), .B2(_1570_ ), .ZN(_1718_ ) );
OAI21_X1 _2614_ ( .A(fanout_net_7 ), .B1(_1573_ ), .B2(_1574_ ), .ZN(_1719_ ) );
NAND2_X1 _2615_ ( .A1(_1718_ ), .A2(_1719_ ), .ZN(_1720_ ) );
NOR2_X1 _2616_ ( .A1(_1576_ ), .A2(fanout_net_7 ), .ZN(_1721_ ) );
MUX2_X1 _2617_ ( .A(_1720_ ), .B(_1721_ ), .S(fanout_net_9 ), .Z(_1722_ ) );
NAND3_X1 _2618_ ( .A1(_1722_ ), .A2(_1676_ ), .A3(_1564_ ), .ZN(_1723_ ) );
NAND2_X1 _2619_ ( .A1(_1581_ ), .A2(_0084_ ), .ZN(_1724_ ) );
BUF_X2 _2620_ ( .A(_1222_ ), .Z(_1725_ ) );
NAND3_X1 _2621_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_1175_ ), .ZN(_1726_ ) );
OAI21_X1 _2622_ ( .A(_1584_ ), .B1(\io_in_a[21] ), .B2(\io_in_b[21] ), .ZN(_1727_ ) );
NAND4_X1 _2623_ ( .A1(_1723_ ), .A2(_1724_ ), .A3(_1726_ ), .A4(_1727_ ), .ZN(_1728_ ) );
NOR4_X1 _2624_ ( .A1(_1687_ ), .A2(_1700_ ), .A3(_1717_ ), .A4(_1728_ ), .ZN(_1729_ ) );
INV_X1 _2625_ ( .A(_1619_ ), .ZN(_1730_ ) );
AND2_X1 _2626_ ( .A1(_1429_ ), .A2(_1423_ ), .ZN(_1731_ ) );
MUX2_X2 _2627_ ( .A(_1731_ ), .B(_1431_ ), .S(fanout_net_5 ), .Z(_1732_ ) );
MUX2_X2 _2628_ ( .A(fanout_net_2 ), .B(_1732_ ), .S(_1611_ ), .Z(_1733_ ) );
OAI211_X1 _2629_ ( .A(fanout_net_12 ), .B(_1602_ ), .C1(_1733_ ), .C2(fanout_net_9 ), .ZN(_1734_ ) );
OAI211_X1 _2630_ ( .A(fanout_net_5 ), .B(_1442_ ), .C1(_1402_ ), .C2(fanout_net_2 ), .ZN(_1735_ ) );
OAI211_X1 _2631_ ( .A(_1275_ ), .B(_1447_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_1736_ ) );
AOI21_X1 _2632_ ( .A(_1240_ ), .B1(_1735_ ), .B2(_1736_ ), .ZN(_1737_ ) );
OAI211_X1 _2633_ ( .A(fanout_net_5 ), .B(_1449_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_1738_ ) );
OAI211_X1 _2634_ ( .A(_1275_ ), .B(_1453_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_1739_ ) );
AOI21_X1 _2635_ ( .A(fanout_net_7 ), .B1(_1738_ ), .B2(_1739_ ), .ZN(_1740_ ) );
OAI21_X1 _2636_ ( .A(_1279_ ), .B1(_1737_ ), .B2(_1740_ ), .ZN(_1741_ ) );
OAI211_X1 _2637_ ( .A(fanout_net_5 ), .B(_1437_ ), .C1(_1296_ ), .C2(fanout_net_2 ), .ZN(_1742_ ) );
OAI211_X1 _2638_ ( .A(_1425_ ), .B(_1440_ ), .C1(_1296_ ), .C2(fanout_net_2 ), .ZN(_1743_ ) );
NAND3_X1 _2639_ ( .A1(_1742_ ), .A2(_1743_ ), .A3(_1211_ ), .ZN(_1744_ ) );
OAI211_X1 _2640_ ( .A(fanout_net_5 ), .B(_1426_ ), .C1(_1296_ ), .C2(fanout_net_2 ), .ZN(_1745_ ) );
OAI211_X1 _2641_ ( .A(_1425_ ), .B(_1435_ ), .C1(_1296_ ), .C2(fanout_net_2 ), .ZN(_1746_ ) );
NAND3_X1 _2642_ ( .A1(_1745_ ), .A2(_1746_ ), .A3(fanout_net_7 ), .ZN(_1747_ ) );
NAND3_X1 _2643_ ( .A1(_1744_ ), .A2(_1747_ ), .A3(fanout_net_9 ), .ZN(_1748_ ) );
NAND2_X1 _2644_ ( .A1(_1741_ ), .A2(_1748_ ), .ZN(_1749_ ) );
NAND2_X1 _2645_ ( .A1(_1749_ ), .A2(_1500_ ), .ZN(_1750_ ) );
AND3_X1 _2646_ ( .A1(_1734_ ), .A2(_1607_ ), .A3(_1750_ ), .ZN(_1751_ ) );
OAI211_X1 _2647_ ( .A(_1683_ ), .B(_1729_ ), .C1(_1730_ ), .C2(_1751_ ), .ZN(\io_out[21] ) );
AND2_X1 _2648_ ( .A1(_1592_ ), .A2(_0073_ ), .ZN(_1752_ ) );
OR3_X1 _2649_ ( .A1(_1752_ ), .A2(_1593_ ), .A3(_1101_ ), .ZN(_1753_ ) );
AOI21_X1 _2650_ ( .A(_1421_ ), .B1(_1355_ ), .B2(fanout_net_2 ), .ZN(_1754_ ) );
INV_X1 _2651_ ( .A(_1754_ ), .ZN(_1755_ ) );
AOI21_X1 _2652_ ( .A(_1601_ ), .B1(_1433_ ), .B2(_1535_ ), .ZN(_1756_ ) );
NAND2_X1 _2653_ ( .A1(_1756_ ), .A2(fanout_net_12 ), .ZN(_1757_ ) );
OAI21_X1 _2654_ ( .A(fanout_net_9 ), .B1(_1439_ ), .B2(_1444_ ), .ZN(_1758_ ) );
OAI21_X1 _2655_ ( .A(_1496_ ), .B1(_1451_ ), .B2(_1457_ ), .ZN(_1759_ ) );
NAND2_X1 _2656_ ( .A1(_1758_ ), .A2(_1759_ ), .ZN(_1760_ ) );
NAND2_X1 _2657_ ( .A1(_1760_ ), .A2(_1676_ ), .ZN(_1761_ ) );
NAND3_X1 _2658_ ( .A1(_1757_ ), .A2(_1421_ ), .A3(_1761_ ), .ZN(_1762_ ) );
AND2_X1 _2659_ ( .A1(_1762_ ), .A2(_1355_ ), .ZN(_1763_ ) );
INV_X1 _2660_ ( .A(_1238_ ), .ZN(_1764_ ) );
AOI21_X1 _2661_ ( .A(_1497_ ), .B1(_1262_ ), .B2(_1267_ ), .ZN(_1765_ ) );
AOI21_X1 _2662_ ( .A(fanout_net_9 ), .B1(_1289_ ), .B2(_1294_ ), .ZN(_1766_ ) );
OAI21_X1 _2663_ ( .A(_1579_ ), .B1(_1765_ ), .B2(_1766_ ), .ZN(_1767_ ) );
AOI211_X1 _2664_ ( .A(fanout_net_7 ), .B(_1257_ ), .C1(_1274_ ), .C2(_1276_ ), .ZN(_1768_ ) );
OAI211_X1 _2665_ ( .A(fanout_net_12 ), .B(_1497_ ), .C1(_1768_ ), .C2(_1273_ ), .ZN(_1769_ ) );
AOI21_X1 _2666_ ( .A(_1764_ ), .B1(_1767_ ), .B2(_1769_ ), .ZN(_1770_ ) );
OAI21_X1 _2667_ ( .A(_1755_ ), .B1(_1763_ ), .B2(_1770_ ), .ZN(_1771_ ) );
AOI21_X1 _2668_ ( .A(_1626_ ), .B1(_1684_ ), .B2(_0073_ ), .ZN(_1772_ ) );
OAI21_X1 _2669_ ( .A(_1772_ ), .B1(_0073_ ), .B2(_1684_ ), .ZN(_1773_ ) );
OAI21_X1 _2670_ ( .A(_1240_ ), .B1(_1329_ ), .B2(_1650_ ), .ZN(_1774_ ) );
OAI21_X1 _2671_ ( .A(fanout_net_7 ), .B1(_1657_ ), .B2(_1658_ ), .ZN(_1775_ ) );
NAND2_X1 _2672_ ( .A1(_1774_ ), .A2(_1775_ ), .ZN(_1776_ ) );
NAND2_X1 _2673_ ( .A1(_1776_ ), .A2(_1321_ ), .ZN(_1777_ ) );
OAI21_X1 _2674_ ( .A(_1327_ ), .B1(_1654_ ), .B2(_1655_ ), .ZN(_1778_ ) );
OAI21_X1 _2675_ ( .A(fanout_net_7 ), .B1(_1668_ ), .B2(_1669_ ), .ZN(_1779_ ) );
NAND2_X1 _2676_ ( .A1(_1778_ ), .A2(_1779_ ), .ZN(_1780_ ) );
NAND2_X1 _2677_ ( .A1(_1780_ ), .A2(fanout_net_9 ), .ZN(_1781_ ) );
AOI21_X1 _2678_ ( .A(_1676_ ), .B1(_1777_ ), .B2(_1781_ ), .ZN(_1782_ ) );
OR3_X1 _2679_ ( .A1(_1300_ ), .A2(_1302_ ), .A3(_1290_ ), .ZN(_1783_ ) );
OR3_X1 _2680_ ( .A1(_1293_ ), .A2(_1299_ ), .A3(fanout_net_7 ), .ZN(_1784_ ) );
AOI21_X1 _2681_ ( .A(fanout_net_9 ), .B1(_1783_ ), .B2(_1784_ ), .ZN(_1785_ ) );
OAI21_X1 _2682_ ( .A(_1240_ ), .B1(_1303_ ), .B2(_1323_ ), .ZN(_1786_ ) );
OAI21_X1 _2683_ ( .A(fanout_net_7 ), .B1(_1325_ ), .B2(_1328_ ), .ZN(_1787_ ) );
AND3_X1 _2684_ ( .A1(_1786_ ), .A2(_1787_ ), .A3(fanout_net_10 ), .ZN(_1788_ ) );
NOR3_X1 _2685_ ( .A1(_1785_ ), .A2(_1788_ ), .A3(fanout_net_12 ), .ZN(_1789_ ) );
OAI21_X1 _2686_ ( .A(_1507_ ), .B1(_1782_ ), .B2(_1789_ ), .ZN(_1790_ ) );
NAND4_X1 _2687_ ( .A1(_1206_ ), .A2(_1510_ ), .A3(\io_in_a[0] ), .A4(fanout_net_10 ), .ZN(_1791_ ) );
OAI21_X1 _2688_ ( .A(_1327_ ), .B1(_1671_ ), .B2(_1672_ ), .ZN(_1792_ ) );
OAI21_X1 _2689_ ( .A(fanout_net_7 ), .B1(_1663_ ), .B2(_1664_ ), .ZN(_1793_ ) );
NAND2_X1 _2690_ ( .A1(_1792_ ), .A2(_1793_ ), .ZN(_1794_ ) );
INV_X1 _2691_ ( .A(_1794_ ), .ZN(_1795_ ) );
OAI21_X1 _2692_ ( .A(_1791_ ), .B1(_1795_ ), .B2(fanout_net_10 ), .ZN(_1796_ ) );
NAND3_X1 _2693_ ( .A1(_1796_ ), .A2(_1677_ ), .A3(_1565_ ), .ZN(_1797_ ) );
OAI21_X1 _2694_ ( .A(_1585_ ), .B1(\io_in_a[20] ), .B2(\io_in_b[20] ), .ZN(_1798_ ) );
AOI22_X1 _2695_ ( .A1(_1176_ ), .A2(_1228_ ), .B1(_1581_ ), .B2(_0073_ ), .ZN(_1799_ ) );
AND4_X1 _2696_ ( .A1(_1790_ ), .A2(_1797_ ), .A3(_1798_ ), .A4(_1799_ ), .ZN(_1800_ ) );
NAND4_X1 _2697_ ( .A1(_1753_ ), .A2(_1771_ ), .A3(_1773_ ), .A4(_1800_ ), .ZN(\io_out[20] ) );
NOR2_X1 _2698_ ( .A1(_1043_ ), .A2(\io_in_b[18] ), .ZN(_1801_ ) );
INV_X1 _2699_ ( .A(_1590_ ), .ZN(_1802_ ) );
OAI21_X1 _2700_ ( .A(_1039_ ), .B1(_1802_ ), .B2(_0234_ ), .ZN(_1803_ ) );
INV_X1 _2701_ ( .A(_0159_ ), .ZN(_1804_ ) );
AOI21_X1 _2702_ ( .A(_1801_ ), .B1(_1803_ ), .B2(_1804_ ), .ZN(_1805_ ) );
AOI21_X1 _2703_ ( .A(_1101_ ), .B1(_1805_ ), .B2(_0191_ ), .ZN(_1806_ ) );
OAI21_X1 _2704_ ( .A(_1806_ ), .B1(_0191_ ), .B2(_1805_ ), .ZN(_1807_ ) );
AOI211_X1 _2705_ ( .A(_1211_ ), .B(_1256_ ), .C1(_1519_ ), .C2(_1521_ ), .ZN(_1808_ ) );
AND4_X1 _2706_ ( .A1(_0589_ ), .A2(_1360_ ), .A3(_1361_ ), .A4(_1696_ ), .ZN(_1809_ ) );
OAI21_X1 _2707_ ( .A(_1209_ ), .B1(_1808_ ), .B2(_1809_ ), .ZN(_1810_ ) );
NAND4_X1 _2708_ ( .A1(_1298_ ), .A2(fanout_net_10 ), .A3(_1318_ ), .A4(_1494_ ), .ZN(_0000_ ) );
AOI21_X1 _2709_ ( .A(_1282_ ), .B1(_1810_ ), .B2(_0000_ ), .ZN(_0001_ ) );
INV_X1 _2710_ ( .A(_0001_ ), .ZN(_0002_ ) );
OAI211_X1 _2711_ ( .A(_1402_ ), .B(fanout_net_7 ), .C1(_1512_ ), .C2(_1508_ ), .ZN(_0003_ ) );
OAI211_X1 _2712_ ( .A(_1402_ ), .B(_1290_ ), .C1(_1514_ ), .C2(_1529_ ), .ZN(_0004_ ) );
AOI21_X1 _2713_ ( .A(_1320_ ), .B1(_0003_ ), .B2(_0004_ ), .ZN(_0005_ ) );
INV_X1 _2714_ ( .A(_0005_ ), .ZN(_0006_ ) );
OAI211_X1 _2715_ ( .A(_1402_ ), .B(fanout_net_7 ), .C1(_1526_ ), .C2(_1531_ ), .ZN(_0007_ ) );
MUX2_X1 _2716_ ( .A(\io_in_a[19] ), .B(\io_in_a[20] ), .S(fanout_net_5 ), .Z(_0008_ ) );
NAND4_X1 _2717_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1290_ ), .A4(_0008_ ), .ZN(_0009_ ) );
AOI21_X1 _2718_ ( .A(fanout_net_10 ), .B1(_0007_ ), .B2(_0009_ ), .ZN(_0010_ ) );
INV_X1 _2719_ ( .A(_0010_ ), .ZN(_0011_ ) );
AOI21_X1 _2720_ ( .A(fanout_net_12 ), .B1(_0006_ ), .B2(_0011_ ), .ZN(_0012_ ) );
INV_X1 _2721_ ( .A(_0012_ ), .ZN(_0013_ ) );
AOI21_X1 _2722_ ( .A(_1688_ ), .B1(_0002_ ), .B2(_0013_ ), .ZN(_0014_ ) );
NOR2_X1 _2723_ ( .A1(_1577_ ), .A2(fanout_net_10 ), .ZN(_0015_ ) );
AND2_X1 _2724_ ( .A1(_0015_ ), .A2(_1214_ ), .ZN(_0016_ ) );
OAI21_X1 _2725_ ( .A(_1218_ ), .B1(_0016_ ), .B2(_1202_ ), .ZN(_0017_ ) );
AOI21_X1 _2726_ ( .A(fanout_net_10 ), .B1(_1548_ ), .B2(_1551_ ), .ZN(_0018_ ) );
AOI21_X1 _2727_ ( .A(_1208_ ), .B1(_1568_ ), .B2(_1571_ ), .ZN(_0019_ ) );
NOR2_X1 _2728_ ( .A1(_0018_ ), .A2(_0019_ ), .ZN(_0020_ ) );
AND3_X1 _2729_ ( .A1(_1556_ ), .A2(fanout_net_10 ), .A3(_1561_ ), .ZN(_0021_ ) );
AOI21_X1 _2730_ ( .A(fanout_net_10 ), .B1(_1539_ ), .B2(_1542_ ), .ZN(_0022_ ) );
OR2_X1 _2731_ ( .A1(_0021_ ), .A2(_0022_ ), .ZN(_0023_ ) );
INV_X1 _2732_ ( .A(_0023_ ), .ZN(_0024_ ) );
MUX2_X1 _2733_ ( .A(_0020_ ), .B(_0024_ ), .S(_1214_ ), .Z(_0025_ ) );
AOI21_X1 _2734_ ( .A(_0017_ ), .B1(_0025_ ), .B2(_1202_ ), .ZN(_0026_ ) );
AND3_X1 _2735_ ( .A1(_1226_ ), .A2(_1222_ ), .A3(_0169_ ), .ZN(_0027_ ) );
AND3_X1 _2736_ ( .A1(_1168_ ), .A2(_1103_ ), .A3(_1231_ ), .ZN(_0028_ ) );
OR4_X1 _2737_ ( .A1(_0014_ ), .A2(_0026_ ), .A3(_0027_ ), .A4(_0028_ ), .ZN(_0029_ ) );
NAND2_X1 _2738_ ( .A1(_1162_ ), .A2(_1166_ ), .ZN(_0031_ ) );
AOI21_X1 _2739_ ( .A(_1804_ ), .B1(_0031_ ), .B2(_1172_ ), .ZN(_0032_ ) );
OR3_X1 _2740_ ( .A1(_0032_ ), .A2(_0191_ ), .A3(_1169_ ), .ZN(_0033_ ) );
OAI21_X1 _2741_ ( .A(_0191_ ), .B1(_0032_ ), .B2(_1169_ ), .ZN(_0034_ ) );
AND3_X1 _2742_ ( .A1(_0033_ ), .A2(_1105_ ), .A3(_0034_ ), .ZN(_0035_ ) );
AOI211_X1 _2743_ ( .A(_0029_ ), .B(_0035_ ), .C1(_0191_ ), .C2(_1582_ ), .ZN(_0036_ ) );
AOI21_X1 _2744_ ( .A(fanout_net_7 ), .B1(_1745_ ), .B2(_1746_ ), .ZN(_0037_ ) );
AOI21_X1 _2745_ ( .A(_0037_ ), .B1(_1732_ ), .B2(fanout_net_7 ), .ZN(_0038_ ) );
AOI21_X1 _2746_ ( .A(_1601_ ), .B1(_0038_ ), .B2(_1496_ ), .ZN(_0039_ ) );
NAND2_X1 _2747_ ( .A1(_0039_ ), .A2(fanout_net_12 ), .ZN(_0040_ ) );
AOI21_X1 _2748_ ( .A(_1212_ ), .B1(_1738_ ), .B2(_1739_ ), .ZN(_0042_ ) );
OAI211_X2 _2749_ ( .A(fanout_net_5 ), .B(_1455_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_0043_ ) );
OAI211_X1 _2750_ ( .A(_1275_ ), .B(_1459_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_0044_ ) );
AOI21_X1 _2751_ ( .A(fanout_net_7 ), .B1(_0043_ ), .B2(_0044_ ), .ZN(_0045_ ) );
OAI21_X1 _2752_ ( .A(_1284_ ), .B1(_0042_ ), .B2(_0045_ ), .ZN(_0046_ ) );
NAND3_X1 _2753_ ( .A1(_1735_ ), .A2(_1736_ ), .A3(_1327_ ), .ZN(_0047_ ) );
NAND3_X1 _2754_ ( .A1(_1742_ ), .A2(_1743_ ), .A3(fanout_net_7 ), .ZN(_0048_ ) );
NAND3_X1 _2755_ ( .A1(_0047_ ), .A2(_0048_ ), .A3(fanout_net_10 ), .ZN(_0049_ ) );
NAND2_X1 _2756_ ( .A1(_0046_ ), .A2(_0049_ ), .ZN(_0050_ ) );
NAND2_X1 _2757_ ( .A1(_0050_ ), .A2(_1283_ ), .ZN(_0051_ ) );
AND3_X1 _2758_ ( .A1(_0040_ ), .A2(_1607_ ), .A3(_0051_ ), .ZN(_0053_ ) );
OAI211_X1 _2759_ ( .A(_1807_ ), .B(_0036_ ), .C1(_1730_ ), .C2(_0053_ ), .ZN(\io_out[19] ) );
AND3_X1 _2760_ ( .A1(_1612_ ), .A2(_1613_ ), .A3(_1320_ ), .ZN(_0054_ ) );
AOI21_X1 _2761_ ( .A(_0054_ ), .B1(_1605_ ), .B2(fanout_net_10 ), .ZN(_0055_ ) );
NOR2_X1 _2762_ ( .A1(_0055_ ), .A2(_1215_ ), .ZN(_0056_ ) );
OAI21_X1 _2763_ ( .A(fanout_net_10 ), .B1(_1608_ ), .B2(_1609_ ), .ZN(_0057_ ) );
AOI21_X1 _2764_ ( .A(_1291_ ), .B1(_1454_ ), .B2(_1456_ ), .ZN(_0058_ ) );
AOI21_X1 _2765_ ( .A(fanout_net_7 ), .B1(_1460_ ), .B2(_1462_ ), .ZN(_0059_ ) );
OAI21_X1 _2766_ ( .A(_1321_ ), .B1(_0058_ ), .B2(_0059_ ), .ZN(_0060_ ) );
AOI21_X1 _2767_ ( .A(fanout_net_12 ), .B1(_0057_ ), .B2(_0060_ ), .ZN(_0061_ ) );
NOR2_X1 _2768_ ( .A1(_0056_ ), .A2(_0061_ ), .ZN(_0063_ ) );
AOI21_X1 _2769_ ( .A(_1356_ ), .B1(_0063_ ), .B2(_1607_ ), .ZN(_0064_ ) );
INV_X1 _2770_ ( .A(_1628_ ), .ZN(_0065_ ) );
INV_X1 _2771_ ( .A(_1629_ ), .ZN(_0066_ ) );
AOI21_X1 _2772_ ( .A(fanout_net_10 ), .B1(_0065_ ), .B2(_0066_ ), .ZN(_0067_ ) );
NOR3_X1 _2773_ ( .A1(_1272_ ), .A2(_1279_ ), .A3(fanout_net_7 ), .ZN(_0068_ ) );
OAI21_X1 _2774_ ( .A(fanout_net_12 ), .B1(_0067_ ), .B2(_0068_ ), .ZN(_0069_ ) );
OAI211_X1 _2775_ ( .A(_1298_ ), .B(fanout_net_7 ), .C1(_1292_ ), .C2(_1293_ ), .ZN(_0070_ ) );
OAI211_X1 _2776_ ( .A(_1298_ ), .B(_1510_ ), .C1(_1299_ ), .C2(_1300_ ), .ZN(_0071_ ) );
NAND2_X1 _2777_ ( .A1(_0070_ ), .A2(_0071_ ), .ZN(_0072_ ) );
NAND2_X1 _2778_ ( .A1(_0072_ ), .A2(_1518_ ), .ZN(_0074_ ) );
AOI21_X1 _2779_ ( .A(_1257_ ), .B1(_1263_ ), .B2(_1265_ ), .ZN(_0075_ ) );
AOI21_X1 _2780_ ( .A(_1633_ ), .B1(fanout_net_7 ), .B2(_0075_ ), .ZN(_0076_ ) );
OAI21_X1 _2781_ ( .A(_0074_ ), .B1(_0076_ ), .B2(_1497_ ), .ZN(_0077_ ) );
NAND2_X1 _2782_ ( .A1(_0077_ ), .A2(_1677_ ), .ZN(_0078_ ) );
AOI21_X1 _2783_ ( .A(_1764_ ), .B1(_0069_ ), .B2(_0078_ ), .ZN(_0079_ ) );
OAI21_X1 _2784_ ( .A(_1755_ ), .B1(_0064_ ), .B2(_0079_ ), .ZN(_0080_ ) );
AOI21_X1 _2785_ ( .A(_1101_ ), .B1(_1803_ ), .B2(_1804_ ), .ZN(_0081_ ) );
OAI21_X1 _2786_ ( .A(_0081_ ), .B1(_1804_ ), .B2(_1803_ ), .ZN(_0082_ ) );
AND3_X1 _2787_ ( .A1(_0031_ ), .A2(_1804_ ), .A3(_1172_ ), .ZN(_0083_ ) );
OR3_X1 _2788_ ( .A1(_0083_ ), .A2(_0032_ ), .A3(_1626_ ), .ZN(_0085_ ) );
AOI21_X1 _2789_ ( .A(fanout_net_10 ), .B1(_1665_ ), .B2(_1666_ ), .ZN(_0086_ ) );
NAND3_X1 _2790_ ( .A1(_1565_ ), .A2(_0086_ ), .A3(_1579_ ), .ZN(_0087_ ) );
OAI21_X1 _2791_ ( .A(_1585_ ), .B1(\io_in_a[18] ), .B2(\io_in_b[18] ), .ZN(_0088_ ) );
AOI22_X1 _2792_ ( .A1(_1169_ ), .A2(_1228_ ), .B1(_1581_ ), .B2(_0159_ ), .ZN(_0089_ ) );
NAND3_X1 _2793_ ( .A1(_0087_ ), .A2(_0088_ ), .A3(_0089_ ), .ZN(_0090_ ) );
NAND2_X1 _2794_ ( .A1(_1674_ ), .A2(fanout_net_10 ), .ZN(_0091_ ) );
NAND3_X1 _2795_ ( .A1(_1656_ ), .A2(_1659_ ), .A3(_1535_ ), .ZN(_0092_ ) );
NAND2_X1 _2796_ ( .A1(_0091_ ), .A2(_0092_ ), .ZN(_0093_ ) );
MUX2_X1 _2797_ ( .A(_1645_ ), .B(_1652_ ), .S(fanout_net_10 ), .Z(_0094_ ) );
MUX2_X1 _2798_ ( .A(_0093_ ), .B(_0094_ ), .S(_1647_ ), .Z(_0096_ ) );
AOI21_X1 _2799_ ( .A(_0090_ ), .B1(_0096_ ), .B2(_1507_ ), .ZN(_0097_ ) );
NAND4_X1 _2800_ ( .A1(_0080_ ), .A2(_0082_ ), .A3(_0085_ ), .A4(_0097_ ), .ZN(\io_out[18] ) );
AND3_X1 _2801_ ( .A1(_1744_ ), .A2(_1747_ ), .A3(_1320_ ), .ZN(_0098_ ) );
AOI21_X2 _2802_ ( .A(_0098_ ), .B1(_1733_ ), .B2(fanout_net_10 ), .ZN(_0099_ ) );
NOR2_X1 _2803_ ( .A1(_0099_ ), .A2(_1215_ ), .ZN(_0100_ ) );
OAI21_X1 _2804_ ( .A(fanout_net_10 ), .B1(_1737_ ), .B2(_1740_ ), .ZN(_0101_ ) );
AOI21_X1 _2805_ ( .A(_1611_ ), .B1(_0043_ ), .B2(_0044_ ), .ZN(_0102_ ) );
OAI211_X1 _2806_ ( .A(fanout_net_5 ), .B(_1461_ ), .C1(_1285_ ), .C2(fanout_net_2 ), .ZN(_0103_ ) );
OAI211_X1 _2807_ ( .A(_1275_ ), .B(_1465_ ), .C1(_1285_ ), .C2(fanout_net_2 ), .ZN(_0104_ ) );
AOI21_X1 _2808_ ( .A(fanout_net_8 ), .B1(_0103_ ), .B2(_0104_ ), .ZN(_0106_ ) );
OAI21_X1 _2809_ ( .A(_1209_ ), .B1(_0102_ ), .B2(_0106_ ), .ZN(_0107_ ) );
AOI21_X1 _2810_ ( .A(fanout_net_12 ), .B1(_0101_ ), .B2(_0107_ ), .ZN(_0108_ ) );
NOR2_X1 _2811_ ( .A1(_0100_ ), .A2(_0108_ ), .ZN(_0109_ ) );
AOI21_X1 _2812_ ( .A(_1356_ ), .B1(_0109_ ), .B2(_1607_ ), .ZN(_0110_ ) );
AOI21_X1 _2813_ ( .A(_1256_ ), .B1(_1519_ ), .B2(_1521_ ), .ZN(_0111_ ) );
AOI21_X1 _2814_ ( .A(_1690_ ), .B1(_0111_ ), .B2(_1211_ ), .ZN(_0112_ ) );
NOR2_X1 _2815_ ( .A1(_0112_ ), .A2(_1535_ ), .ZN(_0113_ ) );
AOI21_X1 _2816_ ( .A(fanout_net_10 ), .B1(_1695_ ), .B2(_1697_ ), .ZN(_0114_ ) );
OAI21_X1 _2817_ ( .A(fanout_net_12 ), .B1(_0113_ ), .B2(_0114_ ), .ZN(_0115_ ) );
AOI21_X1 _2818_ ( .A(_1279_ ), .B1(_1692_ ), .B2(_1693_ ), .ZN(_0117_ ) );
AND4_X1 _2819_ ( .A1(fanout_net_8 ), .A2(_1371_ ), .A3(_1372_ ), .A4(_0008_ ), .ZN(_0118_ ) );
INV_X1 _2820_ ( .A(_0118_ ), .ZN(_0119_ ) );
MUX2_X1 _2821_ ( .A(\io_in_a[17] ), .B(\io_in_a[18] ), .S(fanout_net_5 ), .Z(_0120_ ) );
AND4_X1 _2822_ ( .A1(_1210_ ), .A2(_1371_ ), .A3(_1372_ ), .A4(_0120_ ), .ZN(_0121_ ) );
INV_X1 _2823_ ( .A(_0121_ ), .ZN(_0122_ ) );
AOI21_X1 _2824_ ( .A(fanout_net_10 ), .B1(_0119_ ), .B2(_0122_ ), .ZN(_0123_ ) );
OAI21_X1 _2825_ ( .A(_1283_ ), .B1(_0117_ ), .B2(_0123_ ), .ZN(_0124_ ) );
AOI21_X1 _2826_ ( .A(_1764_ ), .B1(_0115_ ), .B2(_0124_ ), .ZN(_0125_ ) );
OAI21_X1 _2827_ ( .A(_1755_ ), .B1(_0110_ ), .B2(_0125_ ), .ZN(_0126_ ) );
NOR2_X1 _2828_ ( .A1(_1161_ ), .A2(_0289_ ), .ZN(_0128_ ) );
OR3_X1 _2829_ ( .A1(_0128_ ), .A2(_0234_ ), .A3(_0256_ ), .ZN(_0129_ ) );
OAI21_X1 _2830_ ( .A(_0234_ ), .B1(_0128_ ), .B2(_0256_ ), .ZN(_0130_ ) );
NAND3_X1 _2831_ ( .A1(_0129_ ), .A2(_1106_ ), .A3(_0130_ ), .ZN(_0131_ ) );
AOI211_X1 _2832_ ( .A(_1037_ ), .B(_1100_ ), .C1(_1590_ ), .C2(_0245_ ), .ZN(_0132_ ) );
NAND3_X1 _2833_ ( .A1(_1802_ ), .A2(_0234_ ), .A3(_1036_ ), .ZN(_0133_ ) );
NAND2_X1 _2834_ ( .A1(_0132_ ), .A2(_0133_ ), .ZN(_0134_ ) );
AND3_X1 _2835_ ( .A1(_1701_ ), .A2(_1702_ ), .A3(_1351_ ), .ZN(_0135_ ) );
AOI21_X1 _2836_ ( .A(_1351_ ), .B1(_1718_ ), .B2(_1719_ ), .ZN(_0136_ ) );
NOR3_X1 _2837_ ( .A1(_0135_ ), .A2(_1676_ ), .A3(_0136_ ), .ZN(_0137_ ) );
AOI21_X1 _2838_ ( .A(_1320_ ), .B1(_1704_ ), .B2(_1705_ ), .ZN(_0139_ ) );
AND3_X1 _2839_ ( .A1(_1711_ ), .A2(_1712_ ), .A3(_1208_ ), .ZN(_0140_ ) );
OR2_X1 _2840_ ( .A1(_0139_ ), .A2(_0140_ ), .ZN(_0141_ ) );
AOI211_X1 _2841_ ( .A(_1716_ ), .B(_0137_ ), .C1(_1501_ ), .C2(_0141_ ), .ZN(_0142_ ) );
AND4_X1 _2842_ ( .A1(_1579_ ), .A2(_1565_ ), .A3(_1497_ ), .A4(_1721_ ), .ZN(_0143_ ) );
NAND3_X1 _2843_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_0213_ ), .ZN(_0144_ ) );
OAI221_X1 _2844_ ( .A(_0144_ ), .B1(_1234_ ), .B2(_0224_ ), .C1(_1224_ ), .C2(_0245_ ), .ZN(_0145_ ) );
NOR3_X1 _2845_ ( .A1(_0142_ ), .A2(_0143_ ), .A3(_0145_ ), .ZN(_0146_ ) );
NAND4_X1 _2846_ ( .A1(_0126_ ), .A2(_0131_ ), .A3(_0134_ ), .A4(_0146_ ), .ZN(\io_out[17] ) );
NAND3_X1 _2847_ ( .A1(_0931_ ), .A2(_1026_ ), .A3(_0278_ ), .ZN(_0147_ ) );
AND3_X1 _2848_ ( .A1(_1802_ ), .A2(_1487_ ), .A3(_0147_ ), .ZN(_0149_ ) );
AOI21_X1 _2849_ ( .A(_1688_ ), .B1(_1281_ ), .B2(_1306_ ), .ZN(_0150_ ) );
NAND2_X1 _2850_ ( .A1(_1780_ ), .A2(_1284_ ), .ZN(_0151_ ) );
NAND2_X1 _2851_ ( .A1(_1794_ ), .A2(fanout_net_10 ), .ZN(_0152_ ) );
NAND2_X1 _2852_ ( .A1(_0151_ ), .A2(_0152_ ), .ZN(_0153_ ) );
NAND2_X1 _2853_ ( .A1(_0153_ ), .A2(fanout_net_12 ), .ZN(_0154_ ) );
NAND3_X1 _2854_ ( .A1(_1786_ ), .A2(_1787_ ), .A3(_1209_ ), .ZN(_0155_ ) );
OAI21_X1 _2855_ ( .A(_0155_ ), .B1(_1776_ ), .B2(_1351_ ), .ZN(_0156_ ) );
OAI211_X1 _2856_ ( .A(_0154_ ), .B(_1203_ ), .C1(fanout_net_12 ), .C2(_0156_ ), .ZN(_0157_ ) );
INV_X1 _2857_ ( .A(_1218_ ), .ZN(_0158_ ) );
AND2_X1 _2858_ ( .A1(_1213_ ), .A2(_1282_ ), .ZN(_0160_ ) );
INV_X1 _2859_ ( .A(_0160_ ), .ZN(_0161_ ) );
AOI21_X1 _2860_ ( .A(_0158_ ), .B1(_0161_ ), .B2(\io_in_b[4] ), .ZN(_0162_ ) );
AND2_X1 _2861_ ( .A1(_0157_ ), .A2(_0162_ ), .ZN(_0163_ ) );
NAND3_X1 _2862_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_0256_ ), .ZN(_0164_ ) );
OAI221_X1 _2863_ ( .A(_0164_ ), .B1(_1234_ ), .B2(_0267_ ), .C1(_1224_ ), .C2(_0289_ ), .ZN(_0165_ ) );
NOR4_X1 _2864_ ( .A1(_0149_ ), .A2(_0150_ ), .A3(_0163_ ), .A4(_0165_ ), .ZN(_0166_ ) );
AND3_X1 _2865_ ( .A1(_1446_ ), .A2(_1472_ ), .A3(_1421_ ), .ZN(_0167_ ) );
OAI21_X1 _2866_ ( .A(_1106_ ), .B1(_1162_ ), .B2(_0278_ ), .ZN(_0168_ ) );
OAI221_X1 _2867_ ( .A(_0166_ ), .B1(_1730_ ), .B2(_0167_ ), .C1(_0128_ ), .C2(_0168_ ), .ZN(\io_out[16] ) );
INV_X1 _2868_ ( .A(_0697_ ), .ZN(_0170_ ) );
NAND3_X1 _2869_ ( .A1(_1136_ ), .A2(_1140_ ), .A3(_1141_ ), .ZN(_0171_ ) );
AND3_X2 _2870_ ( .A1(_0171_ ), .A2(_1147_ ), .A3(_1152_ ), .ZN(_0172_ ) );
OR4_X4 _2871_ ( .A1(_0170_ ), .A2(_0172_ ), .A3(_0707_ ), .A4(_0718_ ), .ZN(_0173_ ) );
AND2_X2 _2872_ ( .A1(_0173_ ), .A2(_1155_ ), .ZN(_0174_ ) );
OR2_X4 _2873_ ( .A1(_0174_ ), .A2(_0803_ ), .ZN(_0175_ ) );
AND3_X1 _2874_ ( .A1(_0175_ ), .A2(_0782_ ), .A3(_1158_ ), .ZN(_0176_ ) );
AOI21_X4 _2875_ ( .A(_0782_ ), .B1(_0175_ ), .B2(_1158_ ), .ZN(_0177_ ) );
NOR3_X1 _2876_ ( .A1(_0176_ ), .A2(_0177_ ), .A3(_1625_ ), .ZN(_0178_ ) );
OR2_X1 _2877_ ( .A1(_1578_ ), .A2(_1283_ ), .ZN(_0179_ ) );
AND3_X1 _2878_ ( .A1(_0179_ ), .A2(_1506_ ), .A3(_1563_ ), .ZN(_0181_ ) );
NAND3_X1 _2879_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_0750_ ), .ZN(_0182_ ) );
OAI221_X1 _2880_ ( .A(_0182_ ), .B1(_1234_ ), .B2(_0761_ ), .C1(_1224_ ), .C2(_0782_ ), .ZN(_0183_ ) );
INV_X1 _2881_ ( .A(_1239_ ), .ZN(_0184_ ) );
AOI21_X1 _2882_ ( .A(_1809_ ), .B1(_0111_ ), .B2(fanout_net_8 ), .ZN(_0185_ ) );
NOR2_X1 _2883_ ( .A1(_0185_ ), .A2(_1209_ ), .ZN(_0186_ ) );
AOI21_X1 _2884_ ( .A(fanout_net_10 ), .B1(_0003_ ), .B2(_0004_ ), .ZN(_0187_ ) );
OAI21_X1 _2885_ ( .A(fanout_net_12 ), .B1(_0186_ ), .B2(_0187_ ), .ZN(_0188_ ) );
AOI21_X1 _2886_ ( .A(_1284_ ), .B1(_0007_ ), .B2(_0009_ ), .ZN(_0189_ ) );
NAND4_X1 _2887_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(fanout_net_8 ), .A4(_0120_ ), .ZN(_0190_ ) );
MUX2_X1 _2888_ ( .A(\io_in_a[15] ), .B(\io_in_a[16] ), .S(fanout_net_5 ), .Z(_0192_ ) );
NAND4_X1 _2889_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1240_ ), .A4(_0192_ ), .ZN(_0193_ ) );
AOI21_X1 _2890_ ( .A(fanout_net_10 ), .B1(_0190_ ), .B2(_0193_ ), .ZN(_0194_ ) );
OAI21_X1 _2891_ ( .A(_1215_ ), .B1(_0189_ ), .B2(_0194_ ), .ZN(_0195_ ) );
NAND2_X1 _2892_ ( .A1(_0188_ ), .A2(_0195_ ), .ZN(_0196_ ) );
NAND2_X1 _2893_ ( .A1(_0196_ ), .A2(_1203_ ), .ZN(_0197_ ) );
NAND3_X1 _2894_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(fanout_net_2 ), .ZN(_0198_ ) );
NOR3_X1 _2895_ ( .A1(_0198_ ), .A2(\io_in_b[0] ), .A3(fanout_net_8 ), .ZN(_0199_ ) );
NAND4_X1 _2896_ ( .A1(_0199_ ), .A2(\io_in_b[4] ), .A3(_1500_ ), .A4(_1497_ ), .ZN(_0200_ ) );
AOI21_X1 _2897_ ( .A(_0184_ ), .B1(_0197_ ), .B2(_0200_ ), .ZN(_0201_ ) );
NOR4_X1 _2898_ ( .A1(_0178_ ), .A2(_0181_ ), .A3(_0183_ ), .A4(_0201_ ), .ZN(_0203_ ) );
NAND2_X1 _2899_ ( .A1(_0047_ ), .A2(_0048_ ), .ZN(_0204_ ) );
MUX2_X1 _2900_ ( .A(_0204_ ), .B(_0038_ ), .S(fanout_net_10 ), .Z(_0205_ ) );
OAI21_X1 _2901_ ( .A(_1421_ ), .B1(_0205_ ), .B2(_1579_ ), .ZN(_0206_ ) );
OAI21_X1 _2902_ ( .A(fanout_net_10 ), .B1(_0042_ ), .B2(_0045_ ), .ZN(_0207_ ) );
AOI21_X1 _2903_ ( .A(_1212_ ), .B1(_0103_ ), .B2(_0104_ ), .ZN(_0208_ ) );
OAI211_X1 _2904_ ( .A(\io_in_b[0] ), .B(_1467_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_0209_ ) );
OAI211_X1 _2905_ ( .A(_1275_ ), .B(_1362_ ), .C1(_1285_ ), .C2(fanout_net_2 ), .ZN(_0210_ ) );
AOI21_X1 _2906_ ( .A(fanout_net_8 ), .B1(_0209_ ), .B2(_0210_ ), .ZN(_0211_ ) );
OAI21_X1 _2907_ ( .A(_1279_ ), .B1(_0208_ ), .B2(_0211_ ), .ZN(_0212_ ) );
NAND2_X1 _2908_ ( .A1(_0207_ ), .A2(_0212_ ), .ZN(_0214_ ) );
AOI21_X1 _2909_ ( .A(_0206_ ), .B1(_1501_ ), .B2(_0214_ ), .ZN(_0215_ ) );
AND3_X1 _2910_ ( .A1(_0686_ ), .A2(_0867_ ), .A3(_0920_ ), .ZN(_0216_ ) );
NOR2_X1 _2911_ ( .A1(_0216_ ), .A2(_1015_ ), .ZN(_0217_ ) );
NOR2_X1 _2912_ ( .A1(_0217_ ), .A2(_0697_ ), .ZN(_0218_ ) );
AOI21_X1 _2913_ ( .A(_0218_ ), .B1(\io_in_a[12] ), .B2(_1242_ ), .ZN(_0219_ ) );
NOR2_X1 _2914_ ( .A1(_0219_ ), .A2(_0729_ ), .ZN(_0220_ ) );
AOI21_X1 _2915_ ( .A(_0220_ ), .B1(\io_in_a[13] ), .B2(_1019_ ), .ZN(_0221_ ) );
NOR2_X1 _2916_ ( .A1(_0221_ ), .A2(_0793_ ), .ZN(_0222_ ) );
AOI21_X1 _2917_ ( .A(_0222_ ), .B1(\io_in_a[14] ), .B2(_1024_ ), .ZN(_0223_ ) );
AND2_X1 _2918_ ( .A1(_0223_ ), .A2(_0771_ ), .ZN(_0225_ ) );
OAI21_X1 _2919_ ( .A(_1487_ ), .B1(_0223_ ), .B2(_0771_ ), .ZN(_0226_ ) );
OAI221_X1 _2920_ ( .A(_0203_ ), .B1(_1730_ ), .B2(_0215_ ), .C1(_0225_ ), .C2(_0226_ ), .ZN(\io_out[15] ) );
AND2_X1 _2921_ ( .A1(_0221_ ), .A2(_0793_ ), .ZN(_0227_ ) );
OR3_X1 _2922_ ( .A1(_0227_ ), .A2(_0222_ ), .A3(_1101_ ), .ZN(_0228_ ) );
AOI21_X1 _2923_ ( .A(fanout_net_10 ), .B1(_1603_ ), .B2(_1604_ ), .ZN(_0229_ ) );
OAI21_X1 _2924_ ( .A(_1500_ ), .B1(_0229_ ), .B2(_1601_ ), .ZN(_0230_ ) );
NOR2_X1 _2925_ ( .A1(_1214_ ), .A2(fanout_net_2 ), .ZN(_0231_ ) );
INV_X1 _2926_ ( .A(_0231_ ), .ZN(_0232_ ) );
NAND2_X1 _2927_ ( .A1(_0230_ ), .A2(_0232_ ), .ZN(_0233_ ) );
AOI21_X1 _2928_ ( .A(_1359_ ), .B1(_0233_ ), .B2(_1474_ ), .ZN(_0235_ ) );
INV_X1 _2929_ ( .A(_1420_ ), .ZN(_0236_ ) );
BUF_X2 _2930_ ( .A(_0236_ ), .Z(_0237_ ) );
OAI21_X1 _2931_ ( .A(fanout_net_10 ), .B1(_0058_ ), .B2(_0059_ ), .ZN(_0238_ ) );
AOI21_X1 _2932_ ( .A(_1318_ ), .B1(_1466_ ), .B2(_1468_ ), .ZN(_0239_ ) );
AOI21_X1 _2933_ ( .A(fanout_net_8 ), .B1(_1364_ ), .B2(_1366_ ), .ZN(_0240_ ) );
OAI21_X1 _2934_ ( .A(_1518_ ), .B1(_0239_ ), .B2(_0240_ ), .ZN(_0241_ ) );
NAND2_X1 _2935_ ( .A1(_0238_ ), .A2(_0241_ ), .ZN(_0242_ ) );
MUX2_X1 _2936_ ( .A(_1615_ ), .B(_0242_ ), .S(_1647_ ), .Z(_0243_ ) );
OAI21_X1 _2937_ ( .A(_0235_ ), .B1(_0237_ ), .B2(_0243_ ), .ZN(_0244_ ) );
NAND3_X1 _2938_ ( .A1(_1386_ ), .A2(_1387_ ), .A3(\io_in_a[30] ), .ZN(_0246_ ) );
MUX2_X1 _2939_ ( .A(_0198_ ), .B(_0246_ ), .S(_1275_ ), .Z(_0247_ ) );
NOR2_X1 _2940_ ( .A1(_0247_ ), .A2(fanout_net_8 ), .ZN(_0248_ ) );
NAND3_X1 _2941_ ( .A1(_0248_ ), .A2(_1282_ ), .A3(_1321_ ), .ZN(_0249_ ) );
AOI21_X1 _2942_ ( .A(_0184_ ), .B1(_0249_ ), .B2(\io_in_b[4] ), .ZN(_0250_ ) );
AND3_X1 _2943_ ( .A1(_1247_ ), .A2(_1253_ ), .A3(\io_in_a[15] ), .ZN(_0251_ ) );
AND3_X1 _2944_ ( .A1(_1247_ ), .A2(_1253_ ), .A3(\io_in_a[14] ), .ZN(_0252_ ) );
MUX2_X1 _2945_ ( .A(_0251_ ), .B(_0252_ ), .S(_0557_ ), .Z(_0253_ ) );
AND3_X1 _2946_ ( .A1(_1247_ ), .A2(_1253_ ), .A3(\io_in_a[17] ), .ZN(_0254_ ) );
AND3_X1 _2947_ ( .A1(_1247_ ), .A2(_1253_ ), .A3(\io_in_a[16] ), .ZN(_0255_ ) );
MUX2_X1 _2948_ ( .A(_0254_ ), .B(_0255_ ), .S(_0557_ ), .Z(_0257_ ) );
MUX2_X1 _2949_ ( .A(_0253_ ), .B(_0257_ ), .S(fanout_net_8 ), .Z(_0258_ ) );
AND3_X1 _2950_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[21] ), .ZN(_0259_ ) );
AND3_X1 _2951_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[20] ), .ZN(_0260_ ) );
MUX2_X1 _2952_ ( .A(_0259_ ), .B(_0260_ ), .S(_1204_ ), .Z(_0261_ ) );
AND3_X1 _2953_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[19] ), .ZN(_0262_ ) );
AND3_X1 _2954_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[18] ), .ZN(_0263_ ) );
MUX2_X1 _2955_ ( .A(_0262_ ), .B(_0263_ ), .S(_0557_ ), .Z(_0264_ ) );
MUX2_X1 _2956_ ( .A(_0261_ ), .B(_0264_ ), .S(_0589_ ), .Z(_0265_ ) );
MUX2_X1 _2957_ ( .A(_0258_ ), .B(_0265_ ), .S(fanout_net_10 ), .Z(_0266_ ) );
AND3_X1 _2958_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[27] ), .ZN(_0268_ ) );
AND3_X1 _2959_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[26] ), .ZN(_0269_ ) );
MUX2_X1 _2960_ ( .A(_0268_ ), .B(_0269_ ), .S(_1204_ ), .Z(_0270_ ) );
AND3_X1 _2961_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[29] ), .ZN(_0271_ ) );
AND3_X1 _2962_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[28] ), .ZN(_0272_ ) );
MUX2_X1 _2963_ ( .A(_0271_ ), .B(_0272_ ), .S(_0557_ ), .Z(_0273_ ) );
MUX2_X1 _2964_ ( .A(_0270_ ), .B(_0273_ ), .S(fanout_net_8 ), .Z(_0274_ ) );
AND3_X1 _2965_ ( .A1(_1337_ ), .A2(_1339_ ), .A3(\io_in_a[23] ), .ZN(_0275_ ) );
AND3_X1 _2966_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(\io_in_a[22] ), .ZN(_0276_ ) );
MUX2_X1 _2967_ ( .A(_0275_ ), .B(_0276_ ), .S(_1204_ ), .Z(_0277_ ) );
AND3_X1 _2968_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(\io_in_a[25] ), .ZN(_0279_ ) );
AND3_X1 _2969_ ( .A1(_1308_ ), .A2(_1311_ ), .A3(\io_in_a[24] ), .ZN(_0280_ ) );
MUX2_X1 _2970_ ( .A(_0279_ ), .B(_0280_ ), .S(_1204_ ), .Z(_0281_ ) );
MUX2_X1 _2971_ ( .A(_0277_ ), .B(_0281_ ), .S(fanout_net_8 ), .Z(_0282_ ) );
MUX2_X1 _2972_ ( .A(_0274_ ), .B(_0282_ ), .S(_1208_ ), .Z(_0283_ ) );
MUX2_X1 _2973_ ( .A(_0266_ ), .B(_0283_ ), .S(fanout_net_12 ), .Z(_0284_ ) );
OAI21_X1 _2974_ ( .A(_0250_ ), .B1(_0284_ ), .B2(\io_in_b[4] ), .ZN(_0285_ ) );
AND2_X1 _2975_ ( .A1(_1675_ ), .A2(fanout_net_12 ), .ZN(_0286_ ) );
AOI21_X1 _2976_ ( .A(fanout_net_12 ), .B1(_1653_ ), .B2(_1660_ ), .ZN(_0287_ ) );
OAI21_X1 _2977_ ( .A(_1505_ ), .B1(_0286_ ), .B2(_0287_ ), .ZN(_0288_ ) );
NAND3_X1 _2978_ ( .A1(_1226_ ), .A2(_1222_ ), .A3(_1157_ ), .ZN(_0290_ ) );
OAI21_X1 _2979_ ( .A(_1584_ ), .B1(\io_in_a[14] ), .B2(\io_in_b[14] ), .ZN(_0291_ ) );
NAND4_X1 _2980_ ( .A1(_0285_ ), .A2(_0288_ ), .A3(_0290_ ), .A4(_0291_ ), .ZN(_0292_ ) );
AOI21_X1 _2981_ ( .A(_1625_ ), .B1(_0174_ ), .B2(_0803_ ), .ZN(_0293_ ) );
AOI221_X4 _2982_ ( .A(_0292_ ), .B1(_0793_ ), .B2(_1581_ ), .C1(_0175_ ), .C2(_0293_ ), .ZN(_0294_ ) );
NAND3_X1 _2983_ ( .A1(_0228_ ), .A2(_0244_ ), .A3(_0294_ ), .ZN(\io_out[14] ) );
NOR2_X1 _2984_ ( .A1(_1733_ ), .A2(fanout_net_10 ), .ZN(_0295_ ) );
OAI21_X1 _2985_ ( .A(_1283_ ), .B1(_0295_ ), .B2(_1601_ ), .ZN(_0296_ ) );
AND2_X1 _2986_ ( .A1(_0296_ ), .A2(_0232_ ), .ZN(_0297_ ) );
INV_X1 _2987_ ( .A(_1473_ ), .ZN(_0298_ ) );
OAI21_X1 _2988_ ( .A(_1358_ ), .B1(_0297_ ), .B2(_0298_ ), .ZN(_0300_ ) );
AOI21_X1 _2989_ ( .A(_1676_ ), .B1(_1741_ ), .B2(_1748_ ), .ZN(_0301_ ) );
OAI21_X1 _2990_ ( .A(fanout_net_10 ), .B1(_0102_ ), .B2(_0106_ ), .ZN(_0302_ ) );
AOI21_X1 _2991_ ( .A(_1611_ ), .B1(_0209_ ), .B2(_0210_ ), .ZN(_0303_ ) );
OAI211_X2 _2992_ ( .A(\io_in_b[0] ), .B(_1365_ ), .C1(_1285_ ), .C2(fanout_net_2 ), .ZN(_0304_ ) );
OAI211_X1 _2993_ ( .A(_1425_ ), .B(_1369_ ), .C1(_1296_ ), .C2(fanout_net_2 ), .ZN(_0305_ ) );
AOI21_X1 _2994_ ( .A(fanout_net_8 ), .B1(_0304_ ), .B2(_0305_ ), .ZN(_0306_ ) );
OAI21_X1 _2995_ ( .A(_1535_ ), .B1(_0303_ ), .B2(_0306_ ), .ZN(_0307_ ) );
NAND2_X1 _2996_ ( .A1(_0302_ ), .A2(_0307_ ), .ZN(_0308_ ) );
AOI211_X1 _2997_ ( .A(_0237_ ), .B(_0301_ ), .C1(_1501_ ), .C2(_0308_ ), .ZN(_0309_ ) );
OR2_X1 _2998_ ( .A1(_0300_ ), .A2(_0309_ ), .ZN(_0311_ ) );
AND2_X1 _2999_ ( .A1(_0219_ ), .A2(_0729_ ), .ZN(_0312_ ) );
OR3_X1 _3000_ ( .A1(_0312_ ), .A2(_0220_ ), .A3(_1100_ ), .ZN(_0313_ ) );
OR2_X1 _3001_ ( .A1(_0172_ ), .A2(_0170_ ), .ZN(_0314_ ) );
INV_X1 _3002_ ( .A(_1154_ ), .ZN(_0315_ ) );
INV_X1 _3003_ ( .A(_0729_ ), .ZN(_0316_ ) );
AND3_X1 _3004_ ( .A1(_0314_ ), .A2(_0315_ ), .A3(_0316_ ), .ZN(_0317_ ) );
AOI21_X1 _3005_ ( .A(_0316_ ), .B1(_0314_ ), .B2(_0315_ ), .ZN(_0318_ ) );
OR3_X1 _3006_ ( .A1(_0317_ ), .A2(_0318_ ), .A3(_1626_ ), .ZN(_0319_ ) );
NOR3_X1 _3007_ ( .A1(_0112_ ), .A2(fanout_net_13 ), .A3(fanout_net_11 ), .ZN(_0320_ ) );
OAI21_X1 _3008_ ( .A(_1239_ ), .B1(_0320_ ), .B2(_1203_ ), .ZN(_0322_ ) );
NOR2_X1 _3009_ ( .A1(_1694_ ), .A2(_1698_ ), .ZN(_0323_ ) );
NOR2_X1 _3010_ ( .A1(_0118_ ), .A2(_0121_ ), .ZN(_0324_ ) );
AND3_X1 _3011_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[13] ), .ZN(_0325_ ) );
MUX2_X1 _3012_ ( .A(_0252_ ), .B(_0325_ ), .S(_1205_ ), .Z(_0326_ ) );
MUX2_X1 _3013_ ( .A(_0251_ ), .B(_0255_ ), .S(\io_in_b[0] ), .Z(_0327_ ) );
MUX2_X1 _3014_ ( .A(_0326_ ), .B(_0327_ ), .S(fanout_net_8 ), .Z(_0328_ ) );
INV_X1 _3015_ ( .A(_0328_ ), .ZN(_0329_ ) );
MUX2_X1 _3016_ ( .A(_0324_ ), .B(_0329_ ), .S(_1279_ ), .Z(_0330_ ) );
MUX2_X1 _3017_ ( .A(_0323_ ), .B(_0330_ ), .S(_1500_ ), .Z(_0331_ ) );
AOI21_X1 _3018_ ( .A(_0322_ ), .B1(_0331_ ), .B2(_1203_ ), .ZN(_0333_ ) );
OR2_X1 _3019_ ( .A1(_1722_ ), .A2(_1500_ ), .ZN(_0334_ ) );
NAND3_X1 _3020_ ( .A1(_1703_ ), .A2(_1706_ ), .A3(_1676_ ), .ZN(_0335_ ) );
AND3_X1 _3021_ ( .A1(_0334_ ), .A2(_1507_ ), .A3(_0335_ ), .ZN(_0336_ ) );
NAND3_X1 _3022_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_0707_ ), .ZN(_0337_ ) );
OAI221_X1 _3023_ ( .A(_0337_ ), .B1(_1234_ ), .B2(_0718_ ), .C1(_1224_ ), .C2(_0316_ ), .ZN(_0338_ ) );
NOR3_X1 _3024_ ( .A1(_0333_ ), .A2(_0336_ ), .A3(_0338_ ), .ZN(_0339_ ) );
NAND4_X1 _3025_ ( .A1(_0311_ ), .A2(_0313_ ), .A3(_0319_ ), .A4(_0339_ ), .ZN(\io_out[13] ) );
OAI21_X1 _3026_ ( .A(_1105_ ), .B1(_1489_ ), .B2(_1074_ ), .ZN(_0340_ ) );
AOI21_X1 _3027_ ( .A(_0340_ ), .B1(_1074_ ), .B2(_1489_ ), .ZN(_0341_ ) );
AND2_X1 _3028_ ( .A1(_1477_ ), .A2(_1074_ ), .ZN(_0343_ ) );
NOR3_X1 _3029_ ( .A1(_0343_ ), .A2(_1478_ ), .A3(_1100_ ), .ZN(_0344_ ) );
AOI21_X1 _3030_ ( .A(_1730_ ), .B1(_0233_ ), .B2(_1421_ ), .ZN(_0345_ ) );
NOR3_X1 _3031_ ( .A1(_1272_ ), .A2(fanout_net_11 ), .A3(fanout_net_8 ), .ZN(_0346_ ) );
NAND3_X1 _3032_ ( .A1(_0346_ ), .A2(_1216_ ), .A3(_1502_ ), .ZN(_0347_ ) );
OAI21_X1 _3033_ ( .A(_1564_ ), .B1(_0286_ ), .B2(_0287_ ), .ZN(_0348_ ) );
NAND3_X1 _3034_ ( .A1(_1642_ ), .A2(_1646_ ), .A3(fanout_net_13 ), .ZN(_0349_ ) );
OR3_X1 _3035_ ( .A1(_1264_ ), .A2(_1288_ ), .A3(_1611_ ), .ZN(_0350_ ) );
OAI211_X1 _3036_ ( .A(_1263_ ), .B(_1318_ ), .C1(\io_in_b[0] ), .C2(_1065_ ), .ZN(_0351_ ) );
NAND3_X1 _3037_ ( .A1(_0350_ ), .A2(fanout_net_11 ), .A3(_0351_ ), .ZN(_0352_ ) );
OAI211_X1 _3038_ ( .A(_1274_ ), .B(_1510_ ), .C1(\io_in_b[0] ), .C2(_1091_ ), .ZN(_0354_ ) );
NAND2_X1 _3039_ ( .A1(_1276_ ), .A2(_1258_ ), .ZN(_0355_ ) );
OAI211_X1 _3040_ ( .A(_1496_ ), .B(_0354_ ), .C1(_0355_ ), .C2(_1498_ ), .ZN(_0356_ ) );
NAND3_X1 _3041_ ( .A1(_0352_ ), .A2(_1283_ ), .A3(_0356_ ), .ZN(_0357_ ) );
NAND3_X1 _3042_ ( .A1(_0349_ ), .A2(_1506_ ), .A3(_0357_ ), .ZN(_0358_ ) );
OAI21_X1 _3043_ ( .A(_1584_ ), .B1(\io_in_a[30] ), .B2(\io_in_b[30] ), .ZN(_0359_ ) );
NAND2_X1 _3044_ ( .A1(_1223_ ), .A2(_1074_ ), .ZN(_0360_ ) );
NAND3_X1 _3045_ ( .A1(_1226_ ), .A2(_1222_ ), .A3(_1195_ ), .ZN(_0361_ ) );
AND3_X1 _3046_ ( .A1(_0359_ ), .A2(_0360_ ), .A3(_0361_ ), .ZN(_0362_ ) );
NAND4_X1 _3047_ ( .A1(_0347_ ), .A2(_0348_ ), .A3(_0358_ ), .A4(_0362_ ), .ZN(_0363_ ) );
OR4_X1 _3048_ ( .A1(_0341_ ), .A2(_0344_ ), .A3(_0345_ ), .A4(_0363_ ), .ZN(\io_out[30] ) );
NOR3_X1 _3049_ ( .A1(_1278_ ), .A2(fanout_net_13 ), .A3(fanout_net_11 ), .ZN(_0365_ ) );
INV_X1 _3050_ ( .A(_0365_ ), .ZN(_0366_ ) );
AOI21_X1 _3051_ ( .A(_0184_ ), .B1(_0366_ ), .B2(\io_in_b[4] ), .ZN(_0367_ ) );
AOI21_X1 _3052_ ( .A(_1257_ ), .B1(_1258_ ), .B2(_1260_ ), .ZN(_0368_ ) );
MUX2_X1 _3053_ ( .A(_0075_ ), .B(_0368_ ), .S(fanout_net_8 ), .Z(_0369_ ) );
AOI21_X1 _3054_ ( .A(_1766_ ), .B1(_0369_ ), .B2(fanout_net_11 ), .ZN(_0370_ ) );
INV_X1 _3055_ ( .A(_0370_ ), .ZN(_0371_ ) );
AND3_X1 _3056_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(\io_in_a[12] ), .ZN(_0372_ ) );
MUX2_X1 _3057_ ( .A(_0325_ ), .B(_0372_ ), .S(_1205_ ), .Z(_0373_ ) );
MUX2_X1 _3058_ ( .A(_0253_ ), .B(_0373_ ), .S(_1291_ ), .Z(_0375_ ) );
MUX2_X1 _3059_ ( .A(_0264_ ), .B(_0257_ ), .S(_1291_ ), .Z(_0376_ ) );
MUX2_X1 _3060_ ( .A(_0375_ ), .B(_0376_ ), .S(fanout_net_11 ), .Z(_0377_ ) );
MUX2_X1 _3061_ ( .A(_0371_ ), .B(_0377_ ), .S(_1500_ ), .Z(_0378_ ) );
OAI21_X1 _3062_ ( .A(_0367_ ), .B1(_0378_ ), .B2(\io_in_b[4] ), .ZN(_0379_ ) );
NOR3_X1 _3063_ ( .A1(_0216_ ), .A2(_0170_ ), .A3(_1015_ ), .ZN(_0380_ ) );
OR3_X1 _3064_ ( .A1(_0218_ ), .A2(_1100_ ), .A3(_0380_ ), .ZN(_0381_ ) );
AND2_X1 _3065_ ( .A1(_0379_ ), .A2(_0381_ ), .ZN(_0382_ ) );
OAI21_X1 _3066_ ( .A(fanout_net_11 ), .B1(_1463_ ), .B2(_1469_ ), .ZN(_0383_ ) );
OAI21_X1 _3067_ ( .A(_1518_ ), .B1(_1367_ ), .B2(_1375_ ), .ZN(_0384_ ) );
NAND2_X1 _3068_ ( .A1(_0383_ ), .A2(_0384_ ), .ZN(_0386_ ) );
AOI21_X1 _3069_ ( .A(_0237_ ), .B1(_0386_ ), .B2(_1677_ ), .ZN(_0387_ ) );
NAND2_X1 _3070_ ( .A1(_1760_ ), .A2(fanout_net_13 ), .ZN(_0388_ ) );
AOI21_X1 _3071_ ( .A(_1359_ ), .B1(_0387_ ), .B2(_0388_ ), .ZN(_0389_ ) );
NOR2_X1 _3072_ ( .A1(_1756_ ), .A2(fanout_net_13 ), .ZN(_0390_ ) );
NOR2_X1 _3073_ ( .A1(_0390_ ), .A2(_0231_ ), .ZN(_0391_ ) );
OAI21_X1 _3074_ ( .A(_0389_ ), .B1(_0391_ ), .B2(_0298_ ), .ZN(_0392_ ) );
AOI21_X1 _3075_ ( .A(_1626_ ), .B1(_0172_ ), .B2(_0170_ ), .ZN(_0393_ ) );
NAND2_X1 _3076_ ( .A1(_0314_ ), .A2(_0393_ ), .ZN(_0394_ ) );
OAI211_X1 _3077_ ( .A(fanout_net_13 ), .B(_1791_ ), .C1(_1795_ ), .C2(fanout_net_11 ), .ZN(_0395_ ) );
NAND3_X1 _3078_ ( .A1(_1777_ ), .A2(_1781_ ), .A3(_1282_ ), .ZN(_0397_ ) );
NAND3_X1 _3079_ ( .A1(_0395_ ), .A2(_0397_ ), .A3(_1506_ ), .ZN(_0398_ ) );
OAI21_X1 _3080_ ( .A(_1585_ ), .B1(\io_in_a[12] ), .B2(\io_in_b[12] ), .ZN(_0399_ ) );
OAI211_X1 _3081_ ( .A(_0398_ ), .B(_0399_ ), .C1(_0315_ ), .C2(_1229_ ), .ZN(_0400_ ) );
AOI21_X1 _3082_ ( .A(_0400_ ), .B1(_0697_ ), .B2(_1582_ ), .ZN(_0401_ ) );
NAND4_X1 _3083_ ( .A1(_0382_ ), .A2(_0392_ ), .A3(_0394_ ), .A4(_0401_ ), .ZN(\io_out[12] ) );
NOR2_X1 _3084_ ( .A1(_0675_ ), .A2(_0825_ ), .ZN(_0402_ ) );
INV_X1 _3085_ ( .A(_0402_ ), .ZN(_0403_ ) );
OAI21_X1 _3086_ ( .A(_0973_ ), .B1(_0403_ ), .B2(_0857_ ), .ZN(_0404_ ) );
INV_X1 _3087_ ( .A(_0878_ ), .ZN(_0405_ ) );
AND2_X1 _3088_ ( .A1(_0404_ ), .A2(_0405_ ), .ZN(_0407_ ) );
NOR2_X1 _3089_ ( .A1(_1012_ ), .A2(\io_in_b[10] ), .ZN(_0408_ ) );
OR2_X1 _3090_ ( .A1(_0407_ ), .A2(_0408_ ), .ZN(_0409_ ) );
XNOR2_X1 _3091_ ( .A(_0409_ ), .B(_0910_ ), .ZN(_0410_ ) );
NAND2_X1 _3092_ ( .A1(_0410_ ), .A2(_1487_ ), .ZN(_0411_ ) );
NOR2_X1 _3093_ ( .A1(_0039_ ), .A2(fanout_net_13 ), .ZN(_0412_ ) );
OAI21_X1 _3094_ ( .A(_1474_ ), .B1(_0412_ ), .B2(_0231_ ), .ZN(_0413_ ) );
AND2_X1 _3095_ ( .A1(_0413_ ), .A2(_1358_ ), .ZN(_0414_ ) );
OAI21_X1 _3096_ ( .A(fanout_net_11 ), .B1(_0208_ ), .B2(_0211_ ), .ZN(_0415_ ) );
OAI211_X1 _3097_ ( .A(\io_in_b[0] ), .B(_1373_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_0416_ ) );
OAI211_X1 _3098_ ( .A(_1275_ ), .B(_1377_ ), .C1(_1269_ ), .C2(fanout_net_2 ), .ZN(_0418_ ) );
NAND3_X1 _3099_ ( .A1(_0416_ ), .A2(_0418_ ), .A3(_1510_ ), .ZN(_0419_ ) );
NAND3_X1 _3100_ ( .A1(_0304_ ), .A2(_0305_ ), .A3(fanout_net_8 ), .ZN(_0420_ ) );
NAND3_X1 _3101_ ( .A1(_0419_ ), .A2(_0420_ ), .A3(_1518_ ), .ZN(_0421_ ) );
NAND2_X1 _3102_ ( .A1(_0415_ ), .A2(_0421_ ), .ZN(_0422_ ) );
MUX2_X1 _3103_ ( .A(_0422_ ), .B(_0050_ ), .S(fanout_net_13 ), .Z(_0423_ ) );
OAI21_X1 _3104_ ( .A(_0414_ ), .B1(_0237_ ), .B2(_0423_ ), .ZN(_0424_ ) );
AOI21_X1 _3105_ ( .A(_1146_ ), .B1(_1136_ ), .B2(_1140_ ), .ZN(_0425_ ) );
OAI21_X1 _3106_ ( .A(_1150_ ), .B1(_0425_ ), .B2(_0405_ ), .ZN(_0426_ ) );
AOI21_X1 _3107_ ( .A(_1626_ ), .B1(_0426_ ), .B2(_0910_ ), .ZN(_0427_ ) );
OAI21_X1 _3108_ ( .A(_0427_ ), .B1(_0910_ ), .B2(_0426_ ), .ZN(_0429_ ) );
OAI21_X1 _3109_ ( .A(fanout_net_13 ), .B1(_0005_ ), .B2(_0010_ ), .ZN(_0430_ ) );
OAI211_X1 _3110_ ( .A(_1402_ ), .B(fanout_net_8 ), .C1(_1557_ ), .C2(_1555_ ), .ZN(_0431_ ) );
OAI211_X1 _3111_ ( .A(_1402_ ), .B(_1290_ ), .C1(_1546_ ), .C2(_1559_ ), .ZN(_0432_ ) );
AOI21_X1 _3112_ ( .A(fanout_net_11 ), .B1(_0431_ ), .B2(_0432_ ), .ZN(_0433_ ) );
AOI21_X1 _3113_ ( .A(_1321_ ), .B1(_0190_ ), .B2(_0193_ ), .ZN(_0434_ ) );
OAI21_X1 _3114_ ( .A(_1500_ ), .B1(_0433_ ), .B2(_0434_ ), .ZN(_0435_ ) );
NAND2_X1 _3115_ ( .A1(_0430_ ), .A2(_0435_ ), .ZN(_0436_ ) );
NAND2_X1 _3116_ ( .A1(_0436_ ), .A2(_1203_ ), .ZN(_0437_ ) );
OAI21_X1 _3117_ ( .A(_0000_ ), .B1(_0185_ ), .B2(fanout_net_11 ), .ZN(_0438_ ) );
NAND3_X1 _3118_ ( .A1(_0438_ ), .A2(\io_in_b[4] ), .A3(_1579_ ), .ZN(_0440_ ) );
AOI21_X1 _3119_ ( .A(_0184_ ), .B1(_0437_ ), .B2(_0440_ ), .ZN(_0441_ ) );
NAND2_X1 _3120_ ( .A1(_0020_ ), .A2(_1216_ ), .ZN(_0442_ ) );
OAI21_X1 _3121_ ( .A(fanout_net_13 ), .B1(_1577_ ), .B2(fanout_net_11 ), .ZN(_0443_ ) );
AND3_X1 _3122_ ( .A1(_0442_ ), .A2(_1507_ ), .A3(_0443_ ), .ZN(_0444_ ) );
NAND3_X1 _3123_ ( .A1(_0910_ ), .A2(_1104_ ), .A3(_1725_ ), .ZN(_0445_ ) );
OAI221_X1 _3124_ ( .A(_0445_ ), .B1(_1234_ ), .B2(_0899_ ), .C1(_1229_ ), .C2(_1148_ ), .ZN(_0446_ ) );
NOR3_X1 _3125_ ( .A1(_0441_ ), .A2(_0444_ ), .A3(_0446_ ), .ZN(_0447_ ) );
NAND4_X1 _3126_ ( .A1(_0411_ ), .A2(_0424_ ), .A3(_0429_ ), .A4(_0447_ ), .ZN(\io_out[11] ) );
AOI211_X1 _3127_ ( .A(fanout_net_13 ), .B(_0054_ ), .C1(_1605_ ), .C2(fanout_net_11 ), .ZN(_0448_ ) );
NOR2_X1 _3128_ ( .A1(_0448_ ), .A2(_0231_ ), .ZN(_0450_ ) );
OAI21_X1 _3129_ ( .A(_1358_ ), .B1(_0450_ ), .B2(_0298_ ), .ZN(_0451_ ) );
OAI21_X1 _3130_ ( .A(fanout_net_11 ), .B1(_0239_ ), .B2(_0240_ ), .ZN(_0452_ ) );
AOI21_X1 _3131_ ( .A(_1291_ ), .B1(_1370_ ), .B2(_1374_ ), .ZN(_0453_ ) );
AOI21_X1 _3132_ ( .A(fanout_net_8 ), .B1(_1379_ ), .B2(_1381_ ), .ZN(_0454_ ) );
OAI21_X1 _3133_ ( .A(_1321_ ), .B1(_0453_ ), .B2(_0454_ ), .ZN(_0455_ ) );
AOI21_X1 _3134_ ( .A(fanout_net_13 ), .B1(_0452_ ), .B2(_0455_ ), .ZN(_0456_ ) );
AOI21_X1 _3135_ ( .A(_1216_ ), .B1(_0057_ ), .B2(_0060_ ), .ZN(_0457_ ) );
NOR3_X1 _3136_ ( .A1(_0456_ ), .A2(_0457_ ), .A3(_0237_ ), .ZN(_0458_ ) );
OR2_X1 _3137_ ( .A1(_0451_ ), .A2(_0458_ ), .ZN(_0459_ ) );
OAI21_X1 _3138_ ( .A(_1105_ ), .B1(_0425_ ), .B2(_0405_ ), .ZN(_0461_ ) );
AOI21_X1 _3139_ ( .A(_0461_ ), .B1(_0405_ ), .B2(_0425_ ), .ZN(_0462_ ) );
AND3_X1 _3140_ ( .A1(_0878_ ), .A2(_1104_ ), .A3(_1725_ ), .ZN(_0463_ ) );
NAND3_X1 _3141_ ( .A1(_0091_ ), .A2(_0092_ ), .A3(_1500_ ), .ZN(_0464_ ) );
OR2_X1 _3142_ ( .A1(_0086_ ), .A2(_1636_ ), .ZN(_0465_ ) );
NAND3_X1 _3143_ ( .A1(_0464_ ), .A2(_1506_ ), .A3(_0465_ ), .ZN(_0466_ ) );
OAI21_X1 _3144_ ( .A(_1585_ ), .B1(\io_in_a[10] ), .B2(\io_in_b[10] ), .ZN(_0467_ ) );
OAI211_X1 _3145_ ( .A(_0466_ ), .B(_0467_ ), .C1(_1150_ ), .C2(_1229_ ), .ZN(_0468_ ) );
NOR3_X1 _3146_ ( .A1(_0462_ ), .A2(_0463_ ), .A3(_0468_ ), .ZN(_0469_ ) );
AOI21_X1 _3147_ ( .A(_1101_ ), .B1(_0404_ ), .B2(_0405_ ), .ZN(_0470_ ) );
OAI21_X1 _3148_ ( .A(_0470_ ), .B1(_0405_ ), .B2(_0404_ ), .ZN(_0472_ ) );
MUX2_X1 _3149_ ( .A(_0368_ ), .B(_1277_ ), .S(fanout_net_8 ), .Z(_0473_ ) );
AOI21_X1 _3150_ ( .A(_0068_ ), .B1(_0473_ ), .B2(_1518_ ), .ZN(_0474_ ) );
NOR2_X1 _3151_ ( .A1(_0474_ ), .A2(fanout_net_13 ), .ZN(_0475_ ) );
INV_X1 _3152_ ( .A(_0475_ ), .ZN(_0476_ ) );
AOI21_X1 _3153_ ( .A(_0184_ ), .B1(_0476_ ), .B2(\io_in_b[4] ), .ZN(_0477_ ) );
OAI211_X1 _3154_ ( .A(_1298_ ), .B(fanout_net_8 ), .C1(_1302_ ), .C2(_1303_ ), .ZN(_0478_ ) );
OAI211_X1 _3155_ ( .A(_1298_ ), .B(_1498_ ), .C1(_1323_ ), .C2(_1325_ ), .ZN(_0479_ ) );
AOI21_X1 _3156_ ( .A(_1496_ ), .B1(_0478_ ), .B2(_0479_ ), .ZN(_0480_ ) );
OAI211_X1 _3157_ ( .A(_1298_ ), .B(fanout_net_8 ), .C1(_1328_ ), .C2(_1329_ ), .ZN(_0481_ ) );
NAND4_X1 _3158_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1318_ ), .A4(_1316_ ), .ZN(_0483_ ) );
AOI21_X1 _3159_ ( .A(fanout_net_11 ), .B1(_0481_ ), .B2(_0483_ ), .ZN(_0484_ ) );
OR2_X1 _3160_ ( .A1(_0480_ ), .A2(_0484_ ), .ZN(_0485_ ) );
MUX2_X1 _3161_ ( .A(_0485_ ), .B(_0077_ ), .S(fanout_net_13 ), .Z(_0486_ ) );
OAI21_X1 _3162_ ( .A(_0477_ ), .B1(\io_in_b[4] ), .B2(_0486_ ), .ZN(_0487_ ) );
NAND4_X1 _3163_ ( .A1(_0459_ ), .A2(_0469_ ), .A3(_0472_ ), .A4(_0487_ ), .ZN(\io_out[10] ) );
AOI21_X1 _3164_ ( .A(_1144_ ), .B1(_1136_ ), .B2(_0825_ ), .ZN(_0488_ ) );
XNOR2_X1 _3165_ ( .A(_0488_ ), .B(_0857_ ), .ZN(_0489_ ) );
AND2_X1 _3166_ ( .A1(_0489_ ), .A2(_1105_ ), .ZN(_0490_ ) );
NAND2_X1 _3167_ ( .A1(_0099_ ), .A2(_1636_ ), .ZN(_0491_ ) );
NAND2_X1 _3168_ ( .A1(_0491_ ), .A2(_0232_ ), .ZN(_0493_ ) );
AOI21_X1 _3169_ ( .A(_1359_ ), .B1(_0493_ ), .B2(_1474_ ), .ZN(_0494_ ) );
AOI21_X1 _3170_ ( .A(_1282_ ), .B1(_0101_ ), .B2(_0107_ ), .ZN(_0495_ ) );
OAI21_X2 _3171_ ( .A(fanout_net_11 ), .B1(_0303_ ), .B2(_0306_ ), .ZN(_0496_ ) );
OAI211_X2 _3172_ ( .A(\io_in_b[0] ), .B(_1380_ ), .C1(_1402_ ), .C2(fanout_net_2 ), .ZN(_0497_ ) );
OAI211_X1 _3173_ ( .A(_1275_ ), .B(_1384_ ), .C1(_1269_ ), .C2(\io_in_a[31] ), .ZN(_0498_ ) );
NAND3_X1 _3174_ ( .A1(_0497_ ), .A2(_0498_ ), .A3(_1240_ ), .ZN(_0499_ ) );
NAND3_X1 _3175_ ( .A1(_0416_ ), .A2(_0418_ ), .A3(fanout_net_8 ), .ZN(_0500_ ) );
NAND3_X1 _3176_ ( .A1(_0499_ ), .A2(_0500_ ), .A3(_1209_ ), .ZN(_0501_ ) );
AOI21_X1 _3177_ ( .A(fanout_net_13 ), .B1(_0496_ ), .B2(_0501_ ), .ZN(_0502_ ) );
OR4_X2 _3178_ ( .A1(\io_in_b[5] ), .A2(_0495_ ), .A3(_0502_ ), .A4(\io_in_b[4] ), .ZN(_0504_ ) );
AOI221_X2 _3179_ ( .A(_0490_ ), .B1(_0857_ ), .B2(_1581_ ), .C1(_0494_ ), .C2(_0504_ ), .ZN(_0505_ ) );
AOI211_X1 _3180_ ( .A(_0952_ ), .B(_1100_ ), .C1(_0686_ ), .C2(_0867_ ), .ZN(_0506_ ) );
OAI21_X1 _3181_ ( .A(_0857_ ), .B1(_0941_ ), .B2(\io_in_b[8] ), .ZN(_0507_ ) );
OAI21_X1 _3182_ ( .A(_0506_ ), .B1(_0402_ ), .B2(_0507_ ), .ZN(_0508_ ) );
INV_X1 _3183_ ( .A(_0112_ ), .ZN(_0509_ ) );
AOI21_X1 _3184_ ( .A(_0114_ ), .B1(_0509_ ), .B2(fanout_net_11 ), .ZN(_0510_ ) );
OR2_X1 _3185_ ( .A1(_0510_ ), .A2(fanout_net_13 ), .ZN(_0511_ ) );
AOI21_X1 _3186_ ( .A(_0184_ ), .B1(_0511_ ), .B2(\io_in_b[4] ), .ZN(_0512_ ) );
NOR2_X1 _3187_ ( .A1(_0117_ ), .A2(_0123_ ), .ZN(_0513_ ) );
INV_X1 _3188_ ( .A(_0513_ ), .ZN(_0515_ ) );
OAI211_X1 _3189_ ( .A(_1297_ ), .B(fanout_net_8 ), .C1(_1546_ ), .C2(_1559_ ), .ZN(_0516_ ) );
OAI211_X1 _3190_ ( .A(_1297_ ), .B(_1211_ ), .C1(_1549_ ), .C2(_1547_ ), .ZN(_0517_ ) );
AOI21_X1 _3191_ ( .A(fanout_net_11 ), .B1(_0516_ ), .B2(_0517_ ), .ZN(_0518_ ) );
OAI211_X1 _3192_ ( .A(_1297_ ), .B(_1611_ ), .C1(_1557_ ), .C2(_1555_ ), .ZN(_0519_ ) );
NAND4_X1 _3193_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(fanout_net_8 ), .A4(_0192_ ), .ZN(_0520_ ) );
AOI21_X1 _3194_ ( .A(_1496_ ), .B1(_0519_ ), .B2(_0520_ ), .ZN(_0521_ ) );
NOR2_X1 _3195_ ( .A1(_0518_ ), .A2(_0521_ ), .ZN(_0522_ ) );
INV_X1 _3196_ ( .A(_0522_ ), .ZN(_0523_ ) );
MUX2_X1 _3197_ ( .A(_0515_ ), .B(_0523_ ), .S(_1647_ ), .Z(_0524_ ) );
OAI21_X1 _3198_ ( .A(_0512_ ), .B1(\io_in_b[4] ), .B2(_0524_ ), .ZN(_0526_ ) );
NOR2_X1 _3199_ ( .A1(_1234_ ), .A2(_0846_ ), .ZN(_0527_ ) );
OR3_X1 _3200_ ( .A1(_0135_ ), .A2(fanout_net_13 ), .A3(_0136_ ), .ZN(_0528_ ) );
OR3_X1 _3201_ ( .A1(_1576_ ), .A2(fanout_net_11 ), .A3(fanout_net_8 ), .ZN(_0529_ ) );
NAND2_X1 _3202_ ( .A1(_0529_ ), .A2(fanout_net_13 ), .ZN(_0530_ ) );
AND3_X1 _3203_ ( .A1(_0528_ ), .A2(_1506_ ), .A3(_0530_ ), .ZN(_0531_ ) );
AOI211_X1 _3204_ ( .A(_0527_ ), .B(_0531_ ), .C1(_0835_ ), .C2(_1228_ ), .ZN(_0532_ ) );
NAND4_X1 _3205_ ( .A1(_0505_ ), .A2(_0508_ ), .A3(_0526_ ), .A4(_0532_ ), .ZN(\io_out[9] ) );
AOI21_X2 _3206_ ( .A(fanout_net_13 ), .B1(_1434_ ), .B2(_1445_ ), .ZN(_0533_ ) );
OR2_X2 _3207_ ( .A1(_0533_ ), .A2(_0231_ ), .ZN(_0534_ ) );
AOI21_X1 _3208_ ( .A(_1359_ ), .B1(_0534_ ), .B2(_1474_ ), .ZN(_0536_ ) );
OR2_X1 _3209_ ( .A1(_1471_ ), .A2(_1647_ ), .ZN(_0537_ ) );
OAI211_X1 _3210_ ( .A(_0537_ ), .B(_1607_ ), .C1(fanout_net_13 ), .C2(_1392_ ), .ZN(_0538_ ) );
NAND2_X1 _3211_ ( .A1(_0536_ ), .A2(_0538_ ), .ZN(_0539_ ) );
NAND3_X1 _3212_ ( .A1(_0492_ ), .A2(_0664_ ), .A3(_0825_ ), .ZN(_0540_ ) );
NAND3_X1 _3213_ ( .A1(_0403_ ), .A2(_1487_ ), .A3(_0540_ ), .ZN(_0541_ ) );
AOI21_X1 _3214_ ( .A(_1625_ ), .B1(_1136_ ), .B2(_0825_ ), .ZN(_0542_ ) );
OAI21_X1 _3215_ ( .A(_0542_ ), .B1(_0825_ ), .B2(_1136_ ), .ZN(_0543_ ) );
NAND2_X1 _3216_ ( .A1(_0153_ ), .A2(_1636_ ), .ZN(_0544_ ) );
NAND4_X1 _3217_ ( .A1(_1207_ ), .A2(fanout_net_13 ), .A3(_1535_ ), .A4(_1498_ ), .ZN(_0545_ ) );
NAND2_X1 _3218_ ( .A1(_0544_ ), .A2(_0545_ ), .ZN(_0547_ ) );
NAND2_X1 _3219_ ( .A1(_0547_ ), .A2(_1507_ ), .ZN(_0548_ ) );
OAI21_X1 _3220_ ( .A(_1585_ ), .B1(\io_in_a[8] ), .B2(\io_in_b[8] ), .ZN(_0549_ ) );
AOI22_X1 _3221_ ( .A1(_1144_ ), .A2(_1228_ ), .B1(_1582_ ), .B2(_0825_ ), .ZN(_0550_ ) );
AND4_X1 _3222_ ( .A1(_0543_ ), .A2(_0548_ ), .A3(_0549_ ), .A4(_0550_ ), .ZN(_0551_ ) );
OAI211_X1 _3223_ ( .A(\io_in_b[4] ), .B(_1501_ ), .C1(_1268_ ), .C2(_1280_ ), .ZN(_0552_ ) );
OAI21_X1 _3224_ ( .A(fanout_net_13 ), .B1(_1295_ ), .B2(_1305_ ), .ZN(_0553_ ) );
AOI21_X1 _3225_ ( .A(_1518_ ), .B1(_1326_ ), .B2(_1330_ ), .ZN(_0554_ ) );
NAND3_X1 _3226_ ( .A1(_1298_ ), .A2(fanout_net_8 ), .A3(_1316_ ), .ZN(_0555_ ) );
NAND4_X1 _3227_ ( .A1(_1310_ ), .A2(_1313_ ), .A3(_1498_ ), .A4(_1314_ ), .ZN(_0556_ ) );
AOI21_X1 _3228_ ( .A(fanout_net_11 ), .B1(_0555_ ), .B2(_0556_ ), .ZN(_0558_ ) );
OAI21_X1 _3229_ ( .A(_1216_ ), .B1(_0554_ ), .B2(_0558_ ), .ZN(_0559_ ) );
NAND2_X1 _3230_ ( .A1(_0553_ ), .A2(_0559_ ), .ZN(_0560_ ) );
NAND2_X1 _3231_ ( .A1(_0560_ ), .A2(_1203_ ), .ZN(_0561_ ) );
NAND2_X1 _3232_ ( .A1(_0552_ ), .A2(_0561_ ), .ZN(_0562_ ) );
NAND2_X1 _3233_ ( .A1(_0562_ ), .A2(_1239_ ), .ZN(_0563_ ) );
NAND4_X1 _3234_ ( .A1(_0539_ ), .A2(_0541_ ), .A3(_0551_ ), .A4(_0563_ ), .ZN(\io_out[8] ) );
NAND2_X1 _3235_ ( .A1(_0205_ ), .A2(_1283_ ), .ZN(_0564_ ) );
NAND2_X1 _3236_ ( .A1(_0564_ ), .A2(_0232_ ), .ZN(_0565_ ) );
AOI21_X1 _3237_ ( .A(_1359_ ), .B1(_0565_ ), .B2(_1474_ ), .ZN(_0566_ ) );
AOI21_X1 _3238_ ( .A(_0237_ ), .B1(_0214_ ), .B2(fanout_net_13 ), .ZN(_0568_ ) );
OAI211_X1 _3239_ ( .A(\io_in_b[0] ), .B(_1388_ ), .C1(_1363_ ), .C2(\io_in_a[31] ), .ZN(_0569_ ) );
OAI211_X1 _3240_ ( .A(_1259_ ), .B(_1393_ ), .C1(_1378_ ), .C2(\io_in_a[31] ), .ZN(_0570_ ) );
NAND3_X1 _3241_ ( .A1(_0569_ ), .A2(_0570_ ), .A3(_1510_ ), .ZN(_0571_ ) );
NAND3_X1 _3242_ ( .A1(_0497_ ), .A2(_0498_ ), .A3(fanout_net_8 ), .ZN(_0572_ ) );
NAND2_X1 _3243_ ( .A1(_0571_ ), .A2(_0572_ ), .ZN(_0573_ ) );
NAND2_X1 _3244_ ( .A1(_0419_ ), .A2(_0420_ ), .ZN(_0574_ ) );
MUX2_X1 _3245_ ( .A(_0573_ ), .B(_0574_ ), .S(fanout_net_11 ), .Z(_0575_ ) );
OAI21_X1 _3246_ ( .A(_0568_ ), .B1(fanout_net_13 ), .B2(_0575_ ), .ZN(_0576_ ) );
AND2_X1 _3247_ ( .A1(_0566_ ), .A2(_0576_ ), .ZN(_0577_ ) );
AND2_X1 _3248_ ( .A1(_1133_ ), .A2(_0643_ ), .ZN(_0579_ ) );
INV_X1 _3249_ ( .A(_0579_ ), .ZN(_0580_ ) );
AOI21_X1 _3250_ ( .A(_0364_ ), .B1(_0580_ ), .B2(_1118_ ), .ZN(_0581_ ) );
AND2_X1 _3251_ ( .A1(_0581_ ), .A2(_0439_ ), .ZN(_0582_ ) );
INV_X1 _3252_ ( .A(_0582_ ), .ZN(_0583_ ) );
INV_X1 _3253_ ( .A(_1120_ ), .ZN(_0584_ ) );
NAND3_X1 _3254_ ( .A1(_0583_ ), .A2(_0428_ ), .A3(_0584_ ), .ZN(_0585_ ) );
OAI21_X1 _3255_ ( .A(_0460_ ), .B1(_0582_ ), .B2(_1120_ ), .ZN(_0586_ ) );
AOI21_X1 _3256_ ( .A(_1625_ ), .B1(_0585_ ), .B2(_0586_ ), .ZN(_0587_ ) );
AND2_X1 _3257_ ( .A1(_0622_ ), .A2(_0632_ ), .ZN(_0588_ ) );
INV_X1 _3258_ ( .A(_0643_ ), .ZN(_0590_ ) );
INV_X1 _3259_ ( .A(_0374_ ), .ZN(_0591_ ) );
AND3_X1 _3260_ ( .A1(_0588_ ), .A2(_0590_ ), .A3(_0591_ ), .ZN(_0592_ ) );
INV_X1 _3261_ ( .A(_0592_ ), .ZN(_0593_ ) );
AOI21_X1 _3262_ ( .A(_0439_ ), .B1(_0593_ ), .B2(_0417_ ), .ZN(_0594_ ) );
OR3_X1 _3263_ ( .A1(_0594_ ), .A2(_0460_ ), .A3(_0482_ ), .ZN(_0595_ ) );
OAI21_X1 _3264_ ( .A(_0460_ ), .B1(_0594_ ), .B2(_0482_ ), .ZN(_0596_ ) );
AND3_X1 _3265_ ( .A1(_0595_ ), .A2(_1487_ ), .A3(_0596_ ), .ZN(_0597_ ) );
AND2_X1 _3266_ ( .A1(_1238_ ), .A2(_1473_ ), .ZN(_0598_ ) );
INV_X1 _3267_ ( .A(_0598_ ), .ZN(_0599_ ) );
INV_X1 _3268_ ( .A(_0186_ ), .ZN(_0601_ ) );
INV_X1 _3269_ ( .A(_0187_ ), .ZN(_0602_ ) );
AOI21_X1 _3270_ ( .A(fanout_net_13 ), .B1(_0601_ ), .B2(_0602_ ), .ZN(_0603_ ) );
INV_X1 _3271_ ( .A(_0603_ ), .ZN(_0604_ ) );
AND4_X1 _3272_ ( .A1(fanout_net_13 ), .A2(_1495_ ), .A3(_1351_ ), .A4(_1212_ ), .ZN(_0605_ ) );
INV_X1 _3273_ ( .A(_0605_ ), .ZN(_0606_ ) );
AOI21_X1 _3274_ ( .A(_0599_ ), .B1(_0604_ ), .B2(_0606_ ), .ZN(_0607_ ) );
NAND2_X1 _3275_ ( .A1(_0431_ ), .A2(_0432_ ), .ZN(_0608_ ) );
OAI211_X1 _3276_ ( .A(_1255_ ), .B(fanout_net_8 ), .C1(_1549_ ), .C2(_1547_ ), .ZN(_0609_ ) );
OAI211_X1 _3277_ ( .A(_1255_ ), .B(_0589_ ), .C1(_1566_ ), .C2(_1550_ ), .ZN(_0610_ ) );
AND2_X1 _3278_ ( .A1(_0609_ ), .A2(_0610_ ), .ZN(_0612_ ) );
INV_X1 _3279_ ( .A(_0612_ ), .ZN(_0613_ ) );
MUX2_X1 _3280_ ( .A(_0608_ ), .B(_0613_ ), .S(_1320_ ), .Z(_0614_ ) );
OAI21_X1 _3281_ ( .A(_1502_ ), .B1(_0614_ ), .B2(fanout_net_13 ), .ZN(_0615_ ) );
NAND2_X1 _3282_ ( .A1(_0007_ ), .A2(_0009_ ), .ZN(_0616_ ) );
AOI21_X1 _3283_ ( .A(_0194_ ), .B1(_0616_ ), .B2(fanout_net_11 ), .ZN(_0617_ ) );
AOI21_X1 _3284_ ( .A(_0615_ ), .B1(fanout_net_13 ), .B2(_0617_ ), .ZN(_0618_ ) );
NAND3_X1 _3285_ ( .A1(_1578_ ), .A2(_1215_ ), .A3(_1505_ ), .ZN(_0619_ ) );
OAI21_X1 _3286_ ( .A(_1232_ ), .B1(\io_in_a[7] ), .B2(\io_in_b[7] ), .ZN(_0620_ ) );
AOI22_X1 _3287_ ( .A1(_1115_ ), .A2(_1227_ ), .B1(_1223_ ), .B2(_0428_ ), .ZN(_0621_ ) );
NAND3_X1 _3288_ ( .A1(_0619_ ), .A2(_0620_ ), .A3(_0621_ ), .ZN(_0623_ ) );
OR3_X1 _3289_ ( .A1(_0607_ ), .A2(_0618_ ), .A3(_0623_ ), .ZN(_0624_ ) );
OR4_X1 _3290_ ( .A1(_0577_ ), .A2(_0587_ ), .A3(_0597_ ), .A4(_0624_ ), .ZN(\io_out[7] ) );
NAND3_X1 _3291_ ( .A1(_1606_ ), .A2(_1474_ ), .A3(_1616_ ), .ZN(_0625_ ) );
AOI21_X1 _3292_ ( .A(_1216_ ), .B1(_0238_ ), .B2(_0241_ ), .ZN(_0626_ ) );
AOI21_X1 _3293_ ( .A(_1291_ ), .B1(_1385_ ), .B2(_1389_ ), .ZN(_0627_ ) );
AOI21_X1 _3294_ ( .A(fanout_net_8 ), .B1(_1394_ ), .B2(_1396_ ), .ZN(_0628_ ) );
OAI21_X1 _3295_ ( .A(_1518_ ), .B1(_0627_ ), .B2(_0628_ ), .ZN(_0629_ ) );
OAI21_X1 _3296_ ( .A(fanout_net_11 ), .B1(_0453_ ), .B2(_0454_ ), .ZN(_0630_ ) );
AOI21_X1 _3297_ ( .A(fanout_net_13 ), .B1(_0629_ ), .B2(_0630_ ), .ZN(_0631_ ) );
OR3_X1 _3298_ ( .A1(_0626_ ), .A2(_0631_ ), .A3(_0237_ ), .ZN(_0633_ ) );
NAND3_X1 _3299_ ( .A1(_0625_ ), .A2(_1358_ ), .A3(_0633_ ), .ZN(_0634_ ) );
NAND2_X1 _3300_ ( .A1(_1630_ ), .A2(_1634_ ), .ZN(_0635_ ) );
AOI21_X1 _3301_ ( .A(_1637_ ), .B1(_0635_ ), .B2(_1677_ ), .ZN(_0636_ ) );
AOI21_X1 _3302_ ( .A(_0184_ ), .B1(_0636_ ), .B2(\io_in_b[4] ), .ZN(_0637_ ) );
NAND2_X1 _3303_ ( .A1(_0072_ ), .A2(fanout_net_11 ), .ZN(_0638_ ) );
NAND2_X1 _3304_ ( .A1(_0478_ ), .A2(_0479_ ), .ZN(_0639_ ) );
NAND2_X1 _3305_ ( .A1(_0639_ ), .A2(_1497_ ), .ZN(_0640_ ) );
NAND2_X1 _3306_ ( .A1(_0638_ ), .A2(_0640_ ), .ZN(_0641_ ) );
AND2_X1 _3307_ ( .A1(_0481_ ), .A2(_0483_ ), .ZN(_0642_ ) );
INV_X1 _3308_ ( .A(_0642_ ), .ZN(_0644_ ) );
AND3_X1 _3309_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[9] ), .ZN(_0645_ ) );
AND3_X1 _3310_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[8] ), .ZN(_0646_ ) );
MUX2_X1 _3311_ ( .A(_0645_ ), .B(_0646_ ), .S(_1205_ ), .Z(_0647_ ) );
MUX2_X1 _3312_ ( .A(_1335_ ), .B(_0647_ ), .S(fanout_net_8 ), .Z(_0648_ ) );
MUX2_X1 _3313_ ( .A(_0644_ ), .B(_0648_ ), .S(_1535_ ), .Z(_0649_ ) );
MUX2_X1 _3314_ ( .A(_0641_ ), .B(_0649_ ), .S(_1647_ ), .Z(_0650_ ) );
OAI21_X1 _3315_ ( .A(_0637_ ), .B1(_0650_ ), .B2(\io_in_b[4] ), .ZN(_0651_ ) );
OAI21_X1 _3316_ ( .A(_1106_ ), .B1(_0581_ ), .B2(_0439_ ), .ZN(_0652_ ) );
OR2_X1 _3317_ ( .A1(_0582_ ), .A2(_0652_ ), .ZN(_0653_ ) );
NAND3_X1 _3318_ ( .A1(_1675_ ), .A2(_1676_ ), .A3(_1506_ ), .ZN(_0655_ ) );
OAI21_X1 _3319_ ( .A(_1585_ ), .B1(\io_in_a[6] ), .B2(\io_in_b[6] ), .ZN(_0656_ ) );
OAI211_X1 _3320_ ( .A(_0655_ ), .B(_0656_ ), .C1(_0584_ ), .C2(_1229_ ), .ZN(_0657_ ) );
AND3_X1 _3321_ ( .A1(_0593_ ), .A2(_0439_ ), .A3(_0417_ ), .ZN(_0658_ ) );
NOR3_X1 _3322_ ( .A1(_0658_ ), .A2(_0594_ ), .A3(_1100_ ), .ZN(_0659_ ) );
AOI211_X1 _3323_ ( .A(_0657_ ), .B(_0659_ ), .C1(_0439_ ), .C2(_1582_ ), .ZN(_0660_ ) );
NAND4_X1 _3324_ ( .A1(_0634_ ), .A2(_0651_ ), .A3(_0653_ ), .A4(_0660_ ), .ZN(\io_out[6] ) );
AND3_X1 _3325_ ( .A1(_1734_ ), .A2(_1474_ ), .A3(_1750_ ), .ZN(_0661_ ) );
OAI211_X1 _3326_ ( .A(\io_in_b[0] ), .B(_1395_ ), .C1(_1363_ ), .C2(\io_in_a[31] ), .ZN(_0662_ ) );
OAI211_X1 _3327_ ( .A(_1259_ ), .B(_1399_ ), .C1(_1378_ ), .C2(\io_in_a[31] ), .ZN(_0663_ ) );
NAND3_X1 _3328_ ( .A1(_0662_ ), .A2(_0663_ ), .A3(_1291_ ), .ZN(_0665_ ) );
NAND3_X1 _3329_ ( .A1(_0569_ ), .A2(_0570_ ), .A3(\io_in_b[1] ), .ZN(_0666_ ) );
NAND2_X1 _3330_ ( .A1(_0665_ ), .A2(_0666_ ), .ZN(_0667_ ) );
NAND2_X1 _3331_ ( .A1(_0499_ ), .A2(_0500_ ), .ZN(_0668_ ) );
MUX2_X1 _3332_ ( .A(_0667_ ), .B(_0668_ ), .S(fanout_net_11 ), .Z(_0669_ ) );
OAI21_X1 _3333_ ( .A(_1421_ ), .B1(_0669_ ), .B2(fanout_net_13 ), .ZN(_0670_ ) );
AOI21_X1 _3334_ ( .A(_0670_ ), .B1(\io_in_b[3] ), .B2(_0308_ ), .ZN(_0671_ ) );
NOR3_X1 _3335_ ( .A1(_0661_ ), .A2(_1359_ ), .A3(_0671_ ), .ZN(_0672_ ) );
OAI21_X1 _3336_ ( .A(_0374_ ), .B1(_0579_ ), .B2(_1117_ ), .ZN(_0673_ ) );
NAND2_X1 _3337_ ( .A1(_0673_ ), .A2(_1105_ ), .ZN(_0674_ ) );
NOR3_X1 _3338_ ( .A1(_0579_ ), .A2(_1117_ ), .A3(_0374_ ), .ZN(_0676_ ) );
NOR2_X1 _3339_ ( .A1(_0674_ ), .A2(_0676_ ), .ZN(_0677_ ) );
OR3_X1 _3340_ ( .A1(_0592_ ), .A2(_0396_ ), .A3(_1099_ ), .ZN(_0678_ ) );
OAI21_X1 _3341_ ( .A(_0374_ ), .B1(\io_in_b[4] ), .B2(_0385_ ), .ZN(_0679_ ) );
AOI21_X1 _3342_ ( .A(_0679_ ), .B1(_0588_ ), .B2(_0590_ ), .ZN(_0680_ ) );
NOR2_X1 _3343_ ( .A1(_0678_ ), .A2(_0680_ ), .ZN(_0681_ ) );
AND3_X1 _3344_ ( .A1(_1722_ ), .A2(_1215_ ), .A3(_1505_ ), .ZN(_0682_ ) );
NAND3_X1 _3345_ ( .A1(_1226_ ), .A2(_1222_ ), .A3(_0353_ ), .ZN(_0683_ ) );
OAI221_X1 _3346_ ( .A(_0683_ ), .B1(_1234_ ), .B2(_0364_ ), .C1(_1224_ ), .C2(_0591_ ), .ZN(_0684_ ) );
OR3_X1 _3347_ ( .A1(_0681_ ), .A2(_0682_ ), .A3(_0684_ ), .ZN(_0685_ ) );
OAI211_X1 _3348_ ( .A(_1286_ ), .B(\io_in_b[1] ), .C1(_1566_ ), .C2(_1550_ ), .ZN(_0687_ ) );
OAI211_X1 _3349_ ( .A(_1286_ ), .B(_1611_ ), .C1(_1569_ ), .C2(_1567_ ), .ZN(_0688_ ) );
AOI21_X1 _3350_ ( .A(fanout_net_11 ), .B1(_0687_ ), .B2(_0688_ ), .ZN(_0689_ ) );
AOI21_X1 _3351_ ( .A(_1320_ ), .B1(_0516_ ), .B2(_0517_ ), .ZN(_0690_ ) );
OAI21_X1 _3352_ ( .A(_1214_ ), .B1(_0689_ ), .B2(_0690_ ), .ZN(_0691_ ) );
AOI21_X1 _3353_ ( .A(fanout_net_11 ), .B1(_0519_ ), .B2(_0520_ ), .ZN(_0692_ ) );
AOI21_X1 _3354_ ( .A(_1320_ ), .B1(_0119_ ), .B2(_0122_ ), .ZN(_0693_ ) );
OAI21_X1 _3355_ ( .A(\io_in_b[3] ), .B1(_0692_ ), .B2(_0693_ ), .ZN(_0694_ ) );
NAND2_X1 _3356_ ( .A1(_0691_ ), .A2(_0694_ ), .ZN(_0695_ ) );
NOR3_X1 _3357_ ( .A1(_0112_ ), .A2(_1214_ ), .A3(fanout_net_11 ), .ZN(_0696_ ) );
NAND2_X1 _3358_ ( .A1(_1692_ ), .A2(_1693_ ), .ZN(_0698_ ) );
NAND2_X1 _3359_ ( .A1(_0698_ ), .A2(_1320_ ), .ZN(_0699_ ) );
NAND2_X1 _3360_ ( .A1(_1695_ ), .A2(_1697_ ), .ZN(_0700_ ) );
NAND2_X1 _3361_ ( .A1(_0700_ ), .A2(fanout_net_11 ), .ZN(_0701_ ) );
AOI21_X1 _3362_ ( .A(\io_in_b[3] ), .B1(_0699_ ), .B2(_0701_ ), .ZN(_0702_ ) );
NOR2_X1 _3363_ ( .A1(_0696_ ), .A2(_0702_ ), .ZN(_0703_ ) );
INV_X1 _3364_ ( .A(_0703_ ), .ZN(_0704_ ) );
MUX2_X1 _3365_ ( .A(_0695_ ), .B(_0704_ ), .S(\io_in_b[4] ), .Z(_0705_ ) );
AND3_X1 _3366_ ( .A1(_0705_ ), .A2(_0406_ ), .A3(_1238_ ), .ZN(_0706_ ) );
OR4_X1 _3367_ ( .A1(_0672_ ), .A2(_0677_ ), .A3(_0685_ ), .A4(_0706_ ), .ZN(\io_out[5] ) );
NAND3_X1 _3368_ ( .A1(_1757_ ), .A2(_1474_ ), .A3(_1761_ ), .ZN(_0708_ ) );
OAI21_X1 _3369_ ( .A(fanout_net_11 ), .B1(_1382_ ), .B2(_1390_ ), .ZN(_0709_ ) );
OAI211_X1 _3370_ ( .A(_0709_ ), .B(_1647_ ), .C1(_1405_ ), .C2(\io_in_b[2] ), .ZN(_0710_ ) );
OAI21_X1 _3371_ ( .A(_0710_ ), .B1(_1501_ ), .B2(_0386_ ), .ZN(_0711_ ) );
NAND2_X1 _3372_ ( .A1(_0711_ ), .A2(_1607_ ), .ZN(_0712_ ) );
NAND3_X1 _3373_ ( .A1(_0708_ ), .A2(_1358_ ), .A3(_0712_ ), .ZN(_0713_ ) );
AOI21_X1 _3374_ ( .A(_1626_ ), .B1(_1133_ ), .B2(_0643_ ), .ZN(_0714_ ) );
OAI21_X1 _3375_ ( .A(_0714_ ), .B1(_0643_ ), .B2(_1133_ ), .ZN(_0715_ ) );
AOI21_X1 _3376_ ( .A(_1100_ ), .B1(_0588_ ), .B2(_0590_ ), .ZN(_0716_ ) );
OAI21_X1 _3377_ ( .A(_0716_ ), .B1(_0588_ ), .B2(_0590_ ), .ZN(_0717_ ) );
NAND3_X1 _3378_ ( .A1(_1796_ ), .A2(_1677_ ), .A3(_1507_ ), .ZN(_0719_ ) );
OAI21_X1 _3379_ ( .A(_1585_ ), .B1(\io_in_b[4] ), .B2(\io_in_a[4] ), .ZN(_0720_ ) );
AOI22_X1 _3380_ ( .A1(_1117_ ), .A2(_1228_ ), .B1(_1582_ ), .B2(_0643_ ), .ZN(_0721_ ) );
AND4_X1 _3381_ ( .A1(_0717_ ), .A2(_0719_ ), .A3(_0720_ ), .A4(_0721_ ), .ZN(_0722_ ) );
OAI21_X1 _3382_ ( .A(\io_in_b[2] ), .B1(_1261_ ), .B2(_1266_ ), .ZN(_0723_ ) );
NAND2_X1 _3383_ ( .A1(_1289_ ), .A2(_1294_ ), .ZN(_0724_ ) );
NAND2_X1 _3384_ ( .A1(_0724_ ), .A2(_1497_ ), .ZN(_0725_ ) );
AOI21_X1 _3385_ ( .A(\io_in_b[3] ), .B1(_0723_ ), .B2(_0725_ ), .ZN(_0726_ ) );
NOR3_X1 _3386_ ( .A1(_1278_ ), .A2(_1676_ ), .A3(\io_in_b[2] ), .ZN(_0727_ ) );
NOR2_X1 _3387_ ( .A1(_0726_ ), .A2(_0727_ ), .ZN(_0728_ ) );
AOI21_X1 _3388_ ( .A(_0184_ ), .B1(_0728_ ), .B2(\io_in_b[4] ), .ZN(_0730_ ) );
AND3_X1 _3389_ ( .A1(_1338_ ), .A2(_1340_ ), .A3(\io_in_a[11] ), .ZN(_0731_ ) );
AND3_X1 _3390_ ( .A1(_1309_ ), .A2(_1312_ ), .A3(\io_in_a[10] ), .ZN(_0732_ ) );
MUX2_X1 _3391_ ( .A(_0731_ ), .B(_0732_ ), .S(_1205_ ), .Z(_0733_ ) );
MUX2_X1 _3392_ ( .A(_0733_ ), .B(_0647_ ), .S(_1510_ ), .Z(_0734_ ) );
MUX2_X1 _3393_ ( .A(_1343_ ), .B(_0734_ ), .S(\io_in_b[2] ), .Z(_0735_ ) );
MUX2_X1 _3394_ ( .A(_0735_ ), .B(_0377_ ), .S(\io_in_b[3] ), .Z(_0736_ ) );
OAI21_X1 _3395_ ( .A(_0730_ ), .B1(_0736_ ), .B2(\io_in_b[4] ), .ZN(_0737_ ) );
NAND4_X1 _3396_ ( .A1(_0713_ ), .A2(_0715_ ), .A3(_0722_ ), .A4(_0737_ ), .ZN(\io_out[4] ) );
NAND3_X1 _3397_ ( .A1(_0040_ ), .A2(_1473_ ), .A3(_0051_ ), .ZN(_0738_ ) );
NAND2_X1 _3398_ ( .A1(_0738_ ), .A2(_1358_ ), .ZN(_0740_ ) );
AOI21_X1 _3399_ ( .A(_1498_ ), .B1(_0662_ ), .B2(_0663_ ), .ZN(_0741_ ) );
OAI211_X1 _3400_ ( .A(\io_in_b[0] ), .B(_1401_ ), .C1(_1286_ ), .C2(\io_in_a[31] ), .ZN(_0742_ ) );
OAI211_X1 _3401_ ( .A(_1206_ ), .B(_1406_ ), .C1(_1297_ ), .C2(\io_in_a[31] ), .ZN(_0743_ ) );
AOI21_X1 _3402_ ( .A(\io_in_b[1] ), .B1(_0742_ ), .B2(_0743_ ), .ZN(_0744_ ) );
OAI21_X1 _3403_ ( .A(_1535_ ), .B1(_0741_ ), .B2(_0744_ ), .ZN(_0745_ ) );
OAI211_X1 _3404_ ( .A(_0745_ ), .B(_1676_ ), .C1(_1497_ ), .C2(_0573_ ), .ZN(_0746_ ) );
OAI21_X1 _3405_ ( .A(_0746_ ), .B1(_1579_ ), .B2(_0422_ ), .ZN(_0747_ ) );
AOI21_X1 _3406_ ( .A(_0740_ ), .B1(_1607_ ), .B2(_0747_ ), .ZN(_0748_ ) );
OR2_X1 _3407_ ( .A1(_0600_ ), .A2(_0611_ ), .ZN(_0749_ ) );
NAND2_X1 _3408_ ( .A1(_0749_ ), .A2(_0525_ ), .ZN(_0751_ ) );
NOR2_X1 _3409_ ( .A1(_1124_ ), .A2(_1125_ ), .ZN(_0752_ ) );
NOR2_X1 _3410_ ( .A1(_0752_ ), .A2(_1131_ ), .ZN(_0753_ ) );
OAI22_X1 _3411_ ( .A1(_0751_ ), .A2(_1099_ ), .B1(_1625_ ), .B2(_0753_ ), .ZN(_0754_ ) );
AND2_X1 _3412_ ( .A1(_0754_ ), .A2(_1129_ ), .ZN(_0755_ ) );
NAND3_X1 _3413_ ( .A1(_0015_ ), .A2(_1216_ ), .A3(_1506_ ), .ZN(_0756_ ) );
AOI21_X1 _3414_ ( .A(_1233_ ), .B1(_1214_ ), .B2(_0535_ ), .ZN(_0757_ ) );
AOI221_X4 _3415_ ( .A(_0757_ ), .B1(_1128_ ), .B2(_1223_ ), .C1(_1126_ ), .C2(_1227_ ), .ZN(_0758_ ) );
AOI22_X1 _3416_ ( .A1(_0751_ ), .A2(_1098_ ), .B1(_1105_ ), .B2(_0753_ ), .ZN(_0759_ ) );
OAI211_X1 _3417_ ( .A(_0756_ ), .B(_0758_ ), .C1(_0759_ ), .C2(_1129_ ), .ZN(_0760_ ) );
OAI21_X1 _3418_ ( .A(\io_in_b[3] ), .B1(_0433_ ), .B2(_0434_ ), .ZN(_0762_ ) );
OAI21_X1 _3419_ ( .A(_1286_ ), .B1(_1573_ ), .B2(_1570_ ), .ZN(_0763_ ) );
OAI21_X1 _3420_ ( .A(_1286_ ), .B1(_1569_ ), .B2(_1567_ ), .ZN(_0764_ ) );
MUX2_X1 _3421_ ( .A(_0763_ ), .B(_0764_ ), .S(\io_in_b[1] ), .Z(_0765_ ) );
MUX2_X1 _3422_ ( .A(_0612_ ), .B(_0765_ ), .S(_1284_ ), .Z(_0766_ ) );
OAI21_X1 _3423_ ( .A(_0762_ ), .B1(_0766_ ), .B2(\io_in_b[3] ), .ZN(_0767_ ) );
NAND2_X1 _3424_ ( .A1(_0767_ ), .A2(_1503_ ), .ZN(_0768_ ) );
OAI21_X1 _3425_ ( .A(_0598_ ), .B1(_0001_ ), .B2(_0012_ ), .ZN(_0769_ ) );
NAND2_X1 _3426_ ( .A1(_0768_ ), .A2(_0769_ ), .ZN(_0770_ ) );
OR4_X1 _3427_ ( .A1(_0748_ ), .A2(_0755_ ), .A3(_0760_ ), .A4(_0770_ ), .ZN(\io_out[3] ) );
AND2_X1 _3428_ ( .A1(_1073_ ), .A2(_1188_ ), .ZN(_0772_ ) );
NOR2_X1 _3429_ ( .A1(_1084_ ), .A2(\io_in_b[28] ), .ZN(_0773_ ) );
OR3_X1 _3430_ ( .A1(_0772_ ), .A2(_1187_ ), .A3(_0773_ ), .ZN(_0774_ ) );
AOI211_X1 _3431_ ( .A(_1085_ ), .B(_1100_ ), .C1(_1073_ ), .C2(_1080_ ), .ZN(_0775_ ) );
NAND2_X1 _3432_ ( .A1(_0774_ ), .A2(_0775_ ), .ZN(_0776_ ) );
NOR2_X1 _3433_ ( .A1(_1186_ ), .A2(_1188_ ), .ZN(_0777_ ) );
OR3_X1 _3434_ ( .A1(_0777_ ), .A2(_1079_ ), .A3(_1192_ ), .ZN(_0778_ ) );
OAI21_X1 _3435_ ( .A(_1079_ ), .B1(_0777_ ), .B2(_1192_ ), .ZN(_0779_ ) );
NAND3_X1 _3436_ ( .A1(_0778_ ), .A2(_1106_ ), .A3(_0779_ ), .ZN(_0780_ ) );
OAI21_X1 _3437_ ( .A(_1619_ ), .B1(_0297_ ), .B2(_0237_ ), .ZN(_0781_ ) );
NOR2_X1 _3438_ ( .A1(_0112_ ), .A2(\io_in_b[2] ), .ZN(_0783_ ) );
NAND3_X1 _3439_ ( .A1(_0783_ ), .A2(_1677_ ), .A3(_1503_ ), .ZN(_0784_ ) );
OAI211_X1 _3440_ ( .A(_1509_ ), .B(\io_in_b[1] ), .C1(\io_in_b[0] ), .C2(_1063_ ), .ZN(_0785_ ) );
OAI211_X1 _3441_ ( .A(_0785_ ), .B(_1279_ ), .C1(\io_in_b[1] ), .C2(_1523_ ), .ZN(_0786_ ) );
NAND3_X1 _3442_ ( .A1(_1530_ ), .A2(\io_in_b[1] ), .A3(_1532_ ), .ZN(_0787_ ) );
NAND3_X1 _3443_ ( .A1(_1513_ ), .A2(_1611_ ), .A3(_1515_ ), .ZN(_0788_ ) );
NAND3_X1 _3444_ ( .A1(_0787_ ), .A2(_0788_ ), .A3(\io_in_b[2] ), .ZN(_0789_ ) );
NAND3_X1 _3445_ ( .A1(_0786_ ), .A2(_1636_ ), .A3(_0789_ ), .ZN(_0790_ ) );
AND2_X1 _3446_ ( .A1(_0790_ ), .A2(_1506_ ), .ZN(_0791_ ) );
OAI21_X1 _3447_ ( .A(_0791_ ), .B1(_1677_ ), .B2(_1714_ ), .ZN(_0792_ ) );
OAI211_X1 _3448_ ( .A(_1565_ ), .B(_0335_ ), .C1(_1722_ ), .C2(_1647_ ), .ZN(_0794_ ) );
NOR2_X1 _3449_ ( .A1(_1234_ ), .A2(_1078_ ), .ZN(_0795_ ) );
AOI221_X4 _3450_ ( .A(_0795_ ), .B1(_1077_ ), .B2(_1227_ ), .C1(_1079_ ), .C2(_1581_ ), .ZN(_0796_ ) );
AND4_X1 _3451_ ( .A1(_0784_ ), .A2(_0792_ ), .A3(_0794_ ), .A4(_0796_ ), .ZN(_0797_ ) );
NAND4_X1 _3452_ ( .A1(_0776_ ), .A2(_0780_ ), .A3(_0781_ ), .A4(_0797_ ), .ZN(\io_out[29] ) );
NAND2_X1 _3453_ ( .A1(_0600_ ), .A2(_0611_ ), .ZN(_0798_ ) );
NAND3_X1 _3454_ ( .A1(_0749_ ), .A2(_1098_ ), .A3(_0798_ ), .ZN(_0799_ ) );
AOI21_X1 _3455_ ( .A(_1625_ ), .B1(_1124_ ), .B2(_1125_ ), .ZN(_0800_ ) );
OAI21_X1 _3456_ ( .A(_0800_ ), .B1(_1125_ ), .B2(_1124_ ), .ZN(_0801_ ) );
OAI21_X1 _3457_ ( .A(_1584_ ), .B1(\io_in_b[2] ), .B2(\io_in_a[2] ), .ZN(_0802_ ) );
NAND3_X1 _3458_ ( .A1(_0799_ ), .A2(_0801_ ), .A3(_0802_ ), .ZN(_0804_ ) );
AOI21_X1 _3459_ ( .A(_1359_ ), .B1(_0063_ ), .B2(_1474_ ), .ZN(_0805_ ) );
AOI21_X1 _3460_ ( .A(_1282_ ), .B1(_0452_ ), .B2(_0455_ ), .ZN(_0806_ ) );
AOI21_X1 _3461_ ( .A(_1318_ ), .B1(_1400_ ), .B2(_1403_ ), .ZN(_0807_ ) );
AOI21_X1 _3462_ ( .A(\io_in_b[1] ), .B1(_1407_ ), .B2(_1409_ ), .ZN(_0808_ ) );
OAI21_X1 _3463_ ( .A(_1321_ ), .B1(_0807_ ), .B2(_0808_ ), .ZN(_0809_ ) );
OAI21_X1 _3464_ ( .A(\io_in_b[2] ), .B1(_0627_ ), .B2(_0628_ ), .ZN(_0810_ ) );
AOI21_X1 _3465_ ( .A(\io_in_b[3] ), .B1(_0809_ ), .B2(_0810_ ), .ZN(_0811_ ) );
OR3_X1 _3466_ ( .A1(_0806_ ), .A2(_0811_ ), .A3(_0236_ ), .ZN(_0812_ ) );
AOI221_X1 _3467_ ( .A(_0804_ ), .B1(_0611_ ), .B2(_1581_ ), .C1(_0805_ ), .C2(_0812_ ), .ZN(_0813_ ) );
NAND3_X1 _3468_ ( .A1(_1507_ ), .A2(_0086_ ), .A3(_1501_ ), .ZN(_0815_ ) );
NAND3_X1 _3469_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_1131_ ), .ZN(_0816_ ) );
MUX2_X1 _3470_ ( .A(_0248_ ), .B(_0274_ ), .S(_1351_ ), .Z(_0817_ ) );
MUX2_X1 _3471_ ( .A(_0265_ ), .B(_0282_ ), .S(\io_in_b[2] ), .Z(_0818_ ) );
MUX2_X1 _3472_ ( .A(_0817_ ), .B(_0818_ ), .S(_1636_ ), .Z(_0819_ ) );
MUX2_X1 _3473_ ( .A(_1342_ ), .B(_1346_ ), .S(_1611_ ), .Z(_0820_ ) );
MUX2_X1 _3474_ ( .A(_0820_ ), .B(_0648_ ), .S(\io_in_b[2] ), .Z(_0821_ ) );
MUX2_X1 _3475_ ( .A(_0373_ ), .B(_0733_ ), .S(_1240_ ), .Z(_0822_ ) );
MUX2_X1 _3476_ ( .A(_0822_ ), .B(_0258_ ), .S(\io_in_b[2] ), .Z(_0823_ ) );
MUX2_X1 _3477_ ( .A(_0821_ ), .B(_0823_ ), .S(\io_in_b[3] ), .Z(_0824_ ) );
MUX2_X1 _3478_ ( .A(_0819_ ), .B(_0824_ ), .S(_1203_ ), .Z(_0826_ ) );
NAND3_X1 _3479_ ( .A1(_0826_ ), .A2(_0406_ ), .A3(_1238_ ), .ZN(_0827_ ) );
NAND4_X1 _3480_ ( .A1(_0813_ ), .A2(_0815_ ), .A3(_0816_ ), .A4(_0827_ ), .ZN(\io_out[2] ) );
NOR3_X1 _3481_ ( .A1(_0100_ ), .A2(_0298_ ), .A3(_0108_ ), .ZN(_0828_ ) );
OR3_X1 _3482_ ( .A1(_1411_ ), .A2(_1412_ ), .A3(\io_in_a[1] ), .ZN(_0829_ ) );
NAND3_X1 _3483_ ( .A1(_1429_ ), .A2(_1206_ ), .A3(_0829_ ), .ZN(_0830_ ) );
OAI211_X1 _3484_ ( .A(\io_in_b[0] ), .B(_1408_ ), .C1(_1286_ ), .C2(\io_in_a[31] ), .ZN(_0831_ ) );
AOI21_X1 _3485_ ( .A(\io_in_b[1] ), .B1(_0830_ ), .B2(_0831_ ), .ZN(_0832_ ) );
AOI21_X1 _3486_ ( .A(_1318_ ), .B1(_0742_ ), .B2(_0743_ ), .ZN(_0833_ ) );
OAI21_X1 _3487_ ( .A(_1321_ ), .B1(_0832_ ), .B2(_0833_ ), .ZN(_0834_ ) );
OAI211_X1 _3488_ ( .A(_0834_ ), .B(_1215_ ), .C1(_1496_ ), .C2(_0667_ ), .ZN(_0836_ ) );
NAND3_X1 _3489_ ( .A1(_0496_ ), .A2(\io_in_b[3] ), .A3(_0501_ ), .ZN(_0837_ ) );
AOI21_X1 _3490_ ( .A(_0236_ ), .B1(_0836_ ), .B2(_0837_ ), .ZN(_0838_ ) );
OR3_X1 _3491_ ( .A1(_0828_ ), .A2(_1359_ ), .A3(_0838_ ), .ZN(_0839_ ) );
NAND2_X1 _3492_ ( .A1(_1582_ ), .A2(_0546_ ), .ZN(_0840_ ) );
OAI21_X1 _3493_ ( .A(_1585_ ), .B1(\io_in_b[1] ), .B2(\io_in_a[1] ), .ZN(_0841_ ) );
OAI21_X1 _3494_ ( .A(_1098_ ), .B1(_0546_ ), .B2(_0567_ ), .ZN(_0842_ ) );
AOI21_X1 _3495_ ( .A(_0842_ ), .B1(_0546_ ), .B2(_0567_ ), .ZN(_0843_ ) );
XNOR2_X1 _3496_ ( .A(_0546_ ), .B(_1230_ ), .ZN(_0844_ ) );
AOI21_X1 _3497_ ( .A(_0843_ ), .B1(_1106_ ), .B2(_0844_ ), .ZN(_0845_ ) );
AND4_X2 _3498_ ( .A1(_0839_ ), .A2(_0840_ ), .A3(_0841_ ), .A4(_0845_ ), .ZN(_0847_ ) );
OR3_X1 _3499_ ( .A1(_1716_ ), .A2(_0529_ ), .A3(\io_in_b[3] ), .ZN(_0848_ ) );
NAND3_X1 _3500_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_1122_ ), .ZN(_0849_ ) );
NAND2_X1 _3501_ ( .A1(_0115_ ), .A2(_0124_ ), .ZN(_0850_ ) );
MUX2_X1 _3502_ ( .A(_1345_ ), .B(_1347_ ), .S(_1205_ ), .Z(_0851_ ) );
MUX2_X1 _3503_ ( .A(_1341_ ), .B(_1344_ ), .S(_1425_ ), .Z(_0852_ ) );
MUX2_X1 _3504_ ( .A(_0851_ ), .B(_0852_ ), .S(\io_in_b[1] ), .Z(_0853_ ) );
MUX2_X1 _3505_ ( .A(_1334_ ), .B(_1336_ ), .S(_1425_ ), .Z(_0854_ ) );
MUX2_X1 _3506_ ( .A(_1333_ ), .B(_0646_ ), .S(\io_in_b[0] ), .Z(_0855_ ) );
MUX2_X1 _3507_ ( .A(_0854_ ), .B(_0855_ ), .S(\io_in_b[1] ), .Z(_0856_ ) );
MUX2_X1 _3508_ ( .A(_0853_ ), .B(_0856_ ), .S(\io_in_b[2] ), .Z(_0858_ ) );
MUX2_X1 _3509_ ( .A(_0732_ ), .B(_0645_ ), .S(_1425_ ), .Z(_0859_ ) );
MUX2_X1 _3510_ ( .A(_0372_ ), .B(_0731_ ), .S(_1425_ ), .Z(_0860_ ) );
MUX2_X1 _3511_ ( .A(_0859_ ), .B(_0860_ ), .S(\io_in_b[1] ), .Z(_0861_ ) );
MUX2_X1 _3512_ ( .A(_0861_ ), .B(_0328_ ), .S(\io_in_b[2] ), .Z(_0862_ ) );
MUX2_X1 _3513_ ( .A(_0858_ ), .B(_0862_ ), .S(\io_in_b[3] ), .Z(_0863_ ) );
MUX2_X1 _3514_ ( .A(_0850_ ), .B(_0863_ ), .S(_1203_ ), .Z(_0864_ ) );
NAND3_X1 _3515_ ( .A1(_0864_ ), .A2(_0406_ ), .A3(_1238_ ), .ZN(_0865_ ) );
NAND4_X1 _3516_ ( .A1(_0847_ ), .A2(_0848_ ), .A3(_0849_ ), .A4(_0865_ ), .ZN(\io_out[1] ) );
AOI21_X1 _3517_ ( .A(_1101_ ), .B1(_1073_ ), .B2(_1188_ ), .ZN(_0866_ ) );
OAI21_X1 _3518_ ( .A(_0866_ ), .B1(_1188_ ), .B2(_1073_ ), .ZN(_0868_ ) );
OAI21_X1 _3519_ ( .A(_1619_ ), .B1(_0391_ ), .B2(_0237_ ), .ZN(_0869_ ) );
OAI21_X1 _3520_ ( .A(_1105_ ), .B1(_1186_ ), .B2(_1188_ ), .ZN(_0870_ ) );
AOI21_X1 _3521_ ( .A(_0870_ ), .B1(_1188_ ), .B2(_1186_ ), .ZN(_0871_ ) );
NOR2_X1 _3522_ ( .A1(_1278_ ), .A2(\io_in_b[2] ), .ZN(_0872_ ) );
AND3_X1 _3523_ ( .A1(_0872_ ), .A2(_1579_ ), .A3(_1503_ ), .ZN(_0873_ ) );
OAI21_X1 _3524_ ( .A(_1327_ ), .B1(_1264_ ), .B2(_1288_ ), .ZN(_0874_ ) );
OAI21_X1 _3525_ ( .A(\io_in_b[1] ), .B1(_1287_ ), .B2(_1292_ ), .ZN(_0875_ ) );
NAND2_X1 _3526_ ( .A1(_0874_ ), .A2(_0875_ ), .ZN(_0876_ ) );
NAND2_X1 _3527_ ( .A1(_1260_ ), .A2(_1263_ ), .ZN(_0877_ ) );
MUX2_X1 _3528_ ( .A(_0877_ ), .B(_0355_ ), .S(_1212_ ), .Z(_0879_ ) );
MUX2_X1 _3529_ ( .A(_0876_ ), .B(_0879_ ), .S(_1496_ ), .Z(_0880_ ) );
NAND2_X1 _3530_ ( .A1(_0880_ ), .A2(_1647_ ), .ZN(_0881_ ) );
OR3_X1 _3531_ ( .A1(_1785_ ), .A2(_1788_ ), .A3(_1636_ ), .ZN(_0882_ ) );
AOI21_X1 _3532_ ( .A(_1716_ ), .B1(_0881_ ), .B2(_0882_ ), .ZN(_0883_ ) );
AND3_X1 _3533_ ( .A1(_0395_ ), .A2(_0397_ ), .A3(_1564_ ), .ZN(_0884_ ) );
OAI21_X1 _3534_ ( .A(_1584_ ), .B1(\io_in_b[28] ), .B2(\io_in_a[28] ), .ZN(_0885_ ) );
NAND3_X1 _3535_ ( .A1(_1226_ ), .A2(_1222_ ), .A3(_1192_ ), .ZN(_0886_ ) );
OAI211_X1 _3536_ ( .A(_0885_ ), .B(_0886_ ), .C1(_1224_ ), .C2(_1188_ ), .ZN(_0887_ ) );
OR2_X1 _3537_ ( .A1(_0884_ ), .A2(_0887_ ), .ZN(_0888_ ) );
NOR4_X1 _3538_ ( .A1(_0871_ ), .A2(_0873_ ), .A3(_0883_ ), .A4(_0888_ ), .ZN(_0890_ ) );
NAND3_X1 _3539_ ( .A1(_0868_ ), .A2(_0869_ ), .A3(_0890_ ), .ZN(\io_out[28] ) );
INV_X1 _3540_ ( .A(_1060_ ), .ZN(_0891_ ) );
INV_X1 _3541_ ( .A(_1061_ ), .ZN(_0892_ ) );
OAI211_X1 _3542_ ( .A(_0891_ ), .B(_0892_ ), .C1(_1027_ ), .C2(_1051_ ), .ZN(_0893_ ) );
AOI21_X1 _3543_ ( .A(_1055_ ), .B1(_0893_ ), .B2(_1071_ ), .ZN(_0894_ ) );
INV_X1 _3544_ ( .A(_0894_ ), .ZN(_0895_ ) );
OAI21_X1 _3545_ ( .A(_0895_ ), .B1(\io_in_b[26] ), .B2(_1065_ ), .ZN(_0896_ ) );
AND2_X1 _3546_ ( .A1(_0896_ ), .A2(_1054_ ), .ZN(_0897_ ) );
OAI21_X1 _3547_ ( .A(_1487_ ), .B1(_0896_ ), .B2(_1054_ ), .ZN(_0898_ ) );
OR2_X1 _3548_ ( .A1(_0897_ ), .A2(_0898_ ), .ZN(_0900_ ) );
NAND2_X1 _3549_ ( .A1(_1183_ ), .A2(_1184_ ), .ZN(_0901_ ) );
AOI21_X1 _3550_ ( .A(_1056_ ), .B1(_0901_ ), .B2(_1109_ ), .ZN(_0902_ ) );
OR3_X1 _3551_ ( .A1(_0902_ ), .A2(_1053_ ), .A3(_1112_ ), .ZN(_0903_ ) );
OAI21_X1 _3552_ ( .A(_1053_ ), .B1(_0902_ ), .B2(_1112_ ), .ZN(_0904_ ) );
NAND3_X1 _3553_ ( .A1(_0903_ ), .A2(_1106_ ), .A3(_0904_ ), .ZN(_0905_ ) );
OAI21_X1 _3554_ ( .A(_1607_ ), .B1(_0412_ ), .B2(_0231_ ), .ZN(_0906_ ) );
NAND2_X1 _3555_ ( .A1(_0906_ ), .A2(_1619_ ), .ZN(_0907_ ) );
NAND3_X1 _3556_ ( .A1(_0438_ ), .A2(_1677_ ), .A3(_1503_ ), .ZN(_0908_ ) );
AOI21_X1 _3557_ ( .A(_1279_ ), .B1(_1528_ ), .B2(_1533_ ), .ZN(_0909_ ) );
AOI21_X1 _3558_ ( .A(\io_in_b[2] ), .B1(_1511_ ), .B2(_1516_ ), .ZN(_0911_ ) );
OAI21_X1 _3559_ ( .A(_1636_ ), .B1(_0909_ ), .B2(_0911_ ), .ZN(_0912_ ) );
AND2_X1 _3560_ ( .A1(_0912_ ), .A2(_1506_ ), .ZN(_0913_ ) );
OAI21_X1 _3561_ ( .A(_0913_ ), .B1(_1677_ ), .B2(_0023_ ), .ZN(_0914_ ) );
NAND3_X1 _3562_ ( .A1(_0442_ ), .A2(_1565_ ), .A3(_0443_ ), .ZN(_0915_ ) );
AOI22_X1 _3563_ ( .A1(_1111_ ), .A2(_1228_ ), .B1(_1581_ ), .B2(_1053_ ), .ZN(_0916_ ) );
OAI21_X1 _3564_ ( .A(_1584_ ), .B1(\io_in_b[27] ), .B2(\io_in_a[27] ), .ZN(_0917_ ) );
AND2_X1 _3565_ ( .A1(_0916_ ), .A2(_0917_ ), .ZN(_0918_ ) );
AND4_X1 _3566_ ( .A1(_0908_ ), .A2(_0914_ ), .A3(_0915_ ), .A4(_0918_ ), .ZN(_0919_ ) );
NAND4_X1 _3567_ ( .A1(_0900_ ), .A2(_0905_ ), .A3(_0907_ ), .A4(_0919_ ), .ZN(\io_out[27] ) );
AND3_X1 _3568_ ( .A1(_0901_ ), .A2(_1056_ ), .A3(_1109_ ), .ZN(_0921_ ) );
OR3_X1 _3569_ ( .A1(_0921_ ), .A2(_0902_ ), .A3(_1626_ ), .ZN(_0922_ ) );
NAND3_X1 _3570_ ( .A1(_0893_ ), .A2(_1055_ ), .A3(_1071_ ), .ZN(_0923_ ) );
NAND3_X1 _3571_ ( .A1(_0895_ ), .A2(_1487_ ), .A3(_0923_ ), .ZN(_0924_ ) );
OAI21_X1 _3572_ ( .A(_1619_ ), .B1(_0450_ ), .B2(_0237_ ), .ZN(_0925_ ) );
INV_X1 _3573_ ( .A(_0474_ ), .ZN(_0926_ ) );
NAND3_X1 _3574_ ( .A1(_0926_ ), .A2(_1501_ ), .A3(_1503_ ), .ZN(_0927_ ) );
NAND3_X1 _3575_ ( .A1(_0464_ ), .A2(_1565_ ), .A3(_0465_ ), .ZN(_0928_ ) );
OAI21_X1 _3576_ ( .A(_1584_ ), .B1(\io_in_b[26] ), .B2(\io_in_a[26] ), .ZN(_0929_ ) );
NAND3_X1 _3577_ ( .A1(_1484_ ), .A2(_1222_ ), .A3(_1112_ ), .ZN(_0930_ ) );
NAND2_X1 _3578_ ( .A1(_0929_ ), .A2(_0930_ ), .ZN(_0932_ ) );
AND3_X1 _3579_ ( .A1(_0350_ ), .A2(_1351_ ), .A3(_0351_ ), .ZN(_0933_ ) );
AOI21_X1 _3580_ ( .A(_1284_ ), .B1(_1639_ ), .B2(_1640_ ), .ZN(_0934_ ) );
OAI21_X1 _3581_ ( .A(_1636_ ), .B1(_0933_ ), .B2(_0934_ ), .ZN(_0935_ ) );
NAND3_X1 _3582_ ( .A1(_1649_ ), .A2(_1651_ ), .A3(\io_in_b[2] ), .ZN(_0936_ ) );
OAI211_X1 _3583_ ( .A(_0936_ ), .B(\io_in_b[3] ), .C1(_1645_ ), .C2(\io_in_b[2] ), .ZN(_0937_ ) );
AOI21_X1 _3584_ ( .A(_1716_ ), .B1(_0935_ ), .B2(_0937_ ), .ZN(_0938_ ) );
AOI211_X1 _3585_ ( .A(_0932_ ), .B(_0938_ ), .C1(_1055_ ), .C2(_1582_ ), .ZN(_0939_ ) );
AND3_X1 _3586_ ( .A1(_0927_ ), .A2(_0928_ ), .A3(_0939_ ), .ZN(_0940_ ) );
NAND4_X1 _3587_ ( .A1(_0922_ ), .A2(_0924_ ), .A3(_0925_ ), .A4(_0940_ ), .ZN(\io_out[26] ) );
NAND2_X1 _3588_ ( .A1(_1183_ ), .A2(_1061_ ), .ZN(_0942_ ) );
INV_X1 _3589_ ( .A(_1108_ ), .ZN(_0943_ ) );
AND3_X1 _3590_ ( .A1(_0942_ ), .A2(_0891_ ), .A3(_0943_ ), .ZN(_0944_ ) );
AOI21_X1 _3591_ ( .A(_0891_ ), .B1(_0942_ ), .B2(_0943_ ), .ZN(_0945_ ) );
NOR3_X1 _3592_ ( .A1(_0944_ ), .A2(_0945_ ), .A3(_1626_ ), .ZN(_0946_ ) );
OAI21_X1 _3593_ ( .A(_0892_ ), .B1(_1027_ ), .B2(_1051_ ), .ZN(_0947_ ) );
OAI21_X1 _3594_ ( .A(_0947_ ), .B1(\io_in_b[24] ), .B2(_1067_ ), .ZN(_0948_ ) );
OAI21_X1 _3595_ ( .A(_1487_ ), .B1(_0948_ ), .B2(_0891_ ), .ZN(_0949_ ) );
AOI21_X1 _3596_ ( .A(_0949_ ), .B1(_0891_ ), .B2(_0948_ ), .ZN(_0950_ ) );
AOI21_X1 _3597_ ( .A(_1730_ ), .B1(_0493_ ), .B2(_1421_ ), .ZN(_0951_ ) );
INV_X1 _3598_ ( .A(_0510_ ), .ZN(_0953_ ) );
NAND3_X1 _3599_ ( .A1(_0953_ ), .A2(_1647_ ), .A3(_1503_ ), .ZN(_0954_ ) );
NAND3_X1 _3600_ ( .A1(_0528_ ), .A2(_1564_ ), .A3(_0530_ ), .ZN(_0955_ ) );
NAND3_X1 _3601_ ( .A1(_1226_ ), .A2(_1222_ ), .A3(_1058_ ), .ZN(_0956_ ) );
OAI21_X1 _3602_ ( .A(_0956_ ), .B1(_1234_ ), .B2(_1059_ ), .ZN(_0957_ ) );
OR3_X1 _3603_ ( .A1(_0139_ ), .A2(_0140_ ), .A3(_1214_ ), .ZN(_0958_ ) );
AND3_X1 _3604_ ( .A1(_0787_ ), .A2(_0788_ ), .A3(_1320_ ), .ZN(_0959_ ) );
AOI21_X1 _3605_ ( .A(_1209_ ), .B1(_1708_ ), .B2(_1709_ ), .ZN(_0960_ ) );
OAI21_X1 _3606_ ( .A(_1282_ ), .B1(_0959_ ), .B2(_0960_ ), .ZN(_0961_ ) );
AOI21_X1 _3607_ ( .A(_1716_ ), .B1(_0958_ ), .B2(_0961_ ), .ZN(_0962_ ) );
AOI211_X1 _3608_ ( .A(_0957_ ), .B(_0962_ ), .C1(_1060_ ), .C2(_1581_ ), .ZN(_0964_ ) );
NAND3_X1 _3609_ ( .A1(_0954_ ), .A2(_0955_ ), .A3(_0964_ ), .ZN(_0965_ ) );
OR4_X2 _3610_ ( .A1(_0946_ ), .A2(_0950_ ), .A3(_0951_ ), .A4(_0965_ ), .ZN(\io_out[25] ) );
NAND3_X1 _3611_ ( .A1(_1167_ ), .A2(_0892_ ), .A3(_1182_ ), .ZN(_0966_ ) );
AND3_X1 _3612_ ( .A1(_0942_ ), .A2(_1105_ ), .A3(_0966_ ), .ZN(_0967_ ) );
AOI21_X1 _3613_ ( .A(_1730_ ), .B1(_0534_ ), .B2(_1421_ ), .ZN(_0968_ ) );
NAND2_X1 _3614_ ( .A1(_0947_ ), .A2(_1487_ ), .ZN(_0969_ ) );
AOI21_X1 _3615_ ( .A(_0969_ ), .B1(_1061_ ), .B2(_1052_ ), .ZN(_0970_ ) );
AND3_X1 _3616_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(\io_in_a[31] ), .ZN(_0971_ ) );
AND3_X1 _3617_ ( .A1(_1371_ ), .A2(_1372_ ), .A3(\io_in_a[30] ), .ZN(_0972_ ) );
MUX2_X1 _3618_ ( .A(_0971_ ), .B(_0972_ ), .S(_1259_ ), .Z(_0974_ ) );
MUX2_X1 _3619_ ( .A(_0974_ ), .B(_0273_ ), .S(_1212_ ), .Z(_0975_ ) );
MUX2_X1 _3620_ ( .A(_0975_ ), .B(_0369_ ), .S(_1496_ ), .Z(_0976_ ) );
NAND3_X1 _3621_ ( .A1(_0976_ ), .A2(_1216_ ), .A3(_1503_ ), .ZN(_0977_ ) );
NAND2_X1 _3622_ ( .A1(_0547_ ), .A2(_1565_ ), .ZN(_0978_ ) );
NOR2_X1 _3623_ ( .A1(_0156_ ), .A2(_1282_ ), .ZN(_0979_ ) );
NAND2_X1 _3624_ ( .A1(_0876_ ), .A2(_1351_ ), .ZN(_0980_ ) );
NAND3_X1 _3625_ ( .A1(_1783_ ), .A2(_1784_ ), .A3(\io_in_b[2] ), .ZN(_0981_ ) );
AOI21_X1 _3626_ ( .A(\io_in_b[3] ), .B1(_0980_ ), .B2(_0981_ ), .ZN(_0982_ ) );
OAI21_X1 _3627_ ( .A(_1505_ ), .B1(_0979_ ), .B2(_0982_ ), .ZN(_0983_ ) );
OAI21_X1 _3628_ ( .A(_1584_ ), .B1(\io_in_b[24] ), .B2(\io_in_a[24] ), .ZN(_0985_ ) );
AOI22_X1 _3629_ ( .A1(_1108_ ), .A2(_1228_ ), .B1(_1223_ ), .B2(_1061_ ), .ZN(_0986_ ) );
AND3_X1 _3630_ ( .A1(_0983_ ), .A2(_0985_ ), .A3(_0986_ ), .ZN(_0987_ ) );
NAND3_X1 _3631_ ( .A1(_0977_ ), .A2(_0978_ ), .A3(_0987_ ), .ZN(_0988_ ) );
OR4_X2 _3632_ ( .A1(_0967_ ), .A2(_0968_ ), .A3(_0970_ ), .A4(_0988_ ), .ZN(\io_out[24] ) );
OAI21_X2 _3633_ ( .A(_1599_ ), .B1(_1033_ ), .B2(\io_in_b[22] ), .ZN(_0989_ ) );
AOI21_X2 _3634_ ( .A(_1101_ ), .B1(_0989_ ), .B2(_0116_ ), .ZN(_0990_ ) );
OAI21_X1 _3635_ ( .A(_0990_ ), .B1(_0116_ ), .B2(_0989_ ), .ZN(_0991_ ) );
OR3_X1 _3636_ ( .A1(_1624_ ), .A2(_0105_ ), .A3(_1180_ ), .ZN(_0992_ ) );
OAI21_X1 _3637_ ( .A(_0105_ ), .B1(_1624_ ), .B2(_1180_ ), .ZN(_0993_ ) );
NAND3_X1 _3638_ ( .A1(_0992_ ), .A2(_1106_ ), .A3(_0993_ ), .ZN(_0995_ ) );
AND3_X1 _3639_ ( .A1(_1536_ ), .A2(_1501_ ), .A3(_1543_ ), .ZN(_0996_ ) );
AOI21_X1 _3640_ ( .A(_1501_ ), .B1(_1553_ ), .B2(_1562_ ), .ZN(_0997_ ) );
OAI21_X1 _3641_ ( .A(_1507_ ), .B1(_0996_ ), .B2(_0997_ ), .ZN(_0998_ ) );
AOI21_X1 _3642_ ( .A(_1730_ ), .B1(_0565_ ), .B2(_1607_ ), .ZN(_0999_ ) );
OAI21_X1 _3643_ ( .A(_1503_ ), .B1(_0603_ ), .B2(_0605_ ), .ZN(_1000_ ) );
NAND3_X1 _3644_ ( .A1(_1578_ ), .A2(_1579_ ), .A3(_1565_ ), .ZN(_1001_ ) );
NAND2_X1 _3645_ ( .A1(_1582_ ), .A2(_0105_ ), .ZN(_1002_ ) );
OAI21_X1 _3646_ ( .A(_1584_ ), .B1(\io_in_b[23] ), .B2(\io_in_a[23] ), .ZN(_1003_ ) );
NAND3_X1 _3647_ ( .A1(_1484_ ), .A2(_1725_ ), .A3(_1179_ ), .ZN(_1004_ ) );
AND2_X1 _3648_ ( .A1(_1003_ ), .A2(_1004_ ), .ZN(_1006_ ) );
NAND4_X1 _3649_ ( .A1(_1000_ ), .A2(_1001_ ), .A3(_1002_ ), .A4(_1006_ ), .ZN(_1007_ ) );
NOR2_X1 _3650_ ( .A1(_0999_ ), .A2(_1007_ ), .ZN(_1008_ ) );
NAND4_X1 _3651_ ( .A1(_0991_ ), .A2(_0995_ ), .A3(_0998_ ), .A4(_1008_ ), .ZN(\io_out[23] ) );
AOI21_X1 _3652_ ( .A(_1626_ ), .B1(_1491_ ), .B2(_1586_ ), .ZN(_1009_ ) );
OAI21_X1 _3653_ ( .A(_1009_ ), .B1(_0030_ ), .B2(_1491_ ), .ZN(_1010_ ) );
XNOR2_X1 _3654_ ( .A(_1482_ ), .B(_1480_ ), .ZN(_1011_ ) );
OAI21_X1 _3655_ ( .A(_1010_ ), .B1(_1011_ ), .B2(_1101_ ), .ZN(io_overflow ) );
BUF_X8 fanout_buf_1 ( .A(\io_in_a[31] ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(\io_in_a[31] ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\io_in_b[0] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\io_in_b[0] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\io_in_b[0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\io_in_b[1] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\io_in_b[1] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\io_in_b[1] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\io_in_b[2] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\io_in_b[2] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\io_in_b[2] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\io_in_b[3] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\io_in_b[3] ), .Z(fanout_net_13 ) );

endmodule
