//Generate the verilog at 2025-08-31T15:52:45 by iSTA.
module ysyx_25030077_top (
clk,
reset,
ALU_carry,
ALU_overflow,
inst_o
);

input clk ;
input reset ;
output ALU_carry ;
output ALU_overflow ;
output [31:0] inst_o ;

wire clk ;
wire reset ;
wire ALU_carry ;
wire ALU_overflow ;
wire _0000_ ;
wire _0001_ ;
wire _0002_ ;
wire _0003_ ;
wire _0004_ ;
wire _0005_ ;
wire _0006_ ;
wire _0007_ ;
wire _0008_ ;
wire _0009_ ;
wire _0010_ ;
wire _0011_ ;
wire _0012_ ;
wire _0013_ ;
wire _0014_ ;
wire _0015_ ;
wire _0016_ ;
wire _0017_ ;
wire _0018_ ;
wire _0019_ ;
wire _0020_ ;
wire _0021_ ;
wire _0022_ ;
wire _0023_ ;
wire _0024_ ;
wire _0025_ ;
wire _0026_ ;
wire _0027_ ;
wire _0028_ ;
wire _0029_ ;
wire _0030_ ;
wire _0031_ ;
wire _0032_ ;
wire _0033_ ;
wire _0034_ ;
wire _0035_ ;
wire _0036_ ;
wire _0037_ ;
wire _0038_ ;
wire _0039_ ;
wire _0040_ ;
wire _0041_ ;
wire _0042_ ;
wire _0043_ ;
wire _0044_ ;
wire _0045_ ;
wire _0046_ ;
wire _0047_ ;
wire _0048_ ;
wire _0049_ ;
wire _0050_ ;
wire _0051_ ;
wire _0052_ ;
wire _0053_ ;
wire _0054_ ;
wire _0055_ ;
wire _0056_ ;
wire _0057_ ;
wire _0058_ ;
wire _0059_ ;
wire _0060_ ;
wire _0061_ ;
wire _0062_ ;
wire _0063_ ;
wire _0064_ ;
wire _0065_ ;
wire _0066_ ;
wire _0067_ ;
wire _0068_ ;
wire _0069_ ;
wire _0070_ ;
wire _0071_ ;
wire _0072_ ;
wire _0073_ ;
wire _0074_ ;
wire _0075_ ;
wire _0076_ ;
wire _0077_ ;
wire _0078_ ;
wire _0079_ ;
wire _0080_ ;
wire _0081_ ;
wire _0082_ ;
wire _0083_ ;
wire _0084_ ;
wire _0085_ ;
wire _0086_ ;
wire _0087_ ;
wire _0088_ ;
wire _0089_ ;
wire _0090_ ;
wire _0091_ ;
wire _0092_ ;
wire _0093_ ;
wire _0094_ ;
wire _0095_ ;
wire _0096_ ;
wire _0097_ ;
wire _0098_ ;
wire _0099_ ;
wire _0100_ ;
wire _0101_ ;
wire _0102_ ;
wire _0103_ ;
wire _0104_ ;
wire _0105_ ;
wire _0106_ ;
wire _0107_ ;
wire _0108_ ;
wire _0109_ ;
wire _0110_ ;
wire _0111_ ;
wire _0112_ ;
wire _0113_ ;
wire _0114_ ;
wire _0115_ ;
wire _0116_ ;
wire _0117_ ;
wire _0118_ ;
wire _0119_ ;
wire _0120_ ;
wire _0121_ ;
wire _0122_ ;
wire _0123_ ;
wire _0124_ ;
wire _0125_ ;
wire _0126_ ;
wire _0127_ ;
wire _0128_ ;
wire _0129_ ;
wire _0130_ ;
wire _0131_ ;
wire _0132_ ;
wire _0133_ ;
wire _0134_ ;
wire _0135_ ;
wire _0136_ ;
wire _0137_ ;
wire _0138_ ;
wire _0139_ ;
wire _0140_ ;
wire _0141_ ;
wire _0142_ ;
wire _0143_ ;
wire _0144_ ;
wire _0145_ ;
wire _0146_ ;
wire _0147_ ;
wire _0148_ ;
wire _0149_ ;
wire _0150_ ;
wire _0151_ ;
wire _0152_ ;
wire _0153_ ;
wire _0154_ ;
wire _0155_ ;
wire _0156_ ;
wire _0157_ ;
wire _0158_ ;
wire _0159_ ;
wire _0160_ ;
wire _0161_ ;
wire _0162_ ;
wire _0163_ ;
wire _0164_ ;
wire _0165_ ;
wire _0166_ ;
wire _0167_ ;
wire _0168_ ;
wire _0169_ ;
wire _0170_ ;
wire _0171_ ;
wire _0172_ ;
wire _0173_ ;
wire _0174_ ;
wire _0175_ ;
wire _0176_ ;
wire _0177_ ;
wire _0178_ ;
wire _0179_ ;
wire _0180_ ;
wire _0181_ ;
wire _0182_ ;
wire _0183_ ;
wire _0184_ ;
wire _0185_ ;
wire _0186_ ;
wire _0187_ ;
wire _0188_ ;
wire _0189_ ;
wire _0190_ ;
wire _0191_ ;
wire _0192_ ;
wire _0193_ ;
wire _0194_ ;
wire _0195_ ;
wire _0196_ ;
wire _0197_ ;
wire _0198_ ;
wire _0199_ ;
wire _0200_ ;
wire _0201_ ;
wire _0202_ ;
wire _0203_ ;
wire _0204_ ;
wire _0205_ ;
wire _0206_ ;
wire _0207_ ;
wire _0208_ ;
wire _0209_ ;
wire _0210_ ;
wire _0211_ ;
wire _0212_ ;
wire _0213_ ;
wire _0214_ ;
wire _0215_ ;
wire _0216_ ;
wire _0217_ ;
wire _0218_ ;
wire _0219_ ;
wire _0220_ ;
wire _0221_ ;
wire _0222_ ;
wire _0223_ ;
wire _0224_ ;
wire _0225_ ;
wire _0226_ ;
wire _0227_ ;
wire _0228_ ;
wire _0229_ ;
wire _0230_ ;
wire _0231_ ;
wire _0232_ ;
wire _0233_ ;
wire _0234_ ;
wire _0235_ ;
wire _0236_ ;
wire _0237_ ;
wire _0238_ ;
wire _0239_ ;
wire _0240_ ;
wire _0241_ ;
wire _0242_ ;
wire _0243_ ;
wire _0244_ ;
wire _0245_ ;
wire _0246_ ;
wire _0247_ ;
wire _0248_ ;
wire _0249_ ;
wire _0250_ ;
wire _0251_ ;
wire _0252_ ;
wire _0253_ ;
wire _0254_ ;
wire _0255_ ;
wire _0256_ ;
wire _0257_ ;
wire _0258_ ;
wire _0259_ ;
wire _0260_ ;
wire _0261_ ;
wire _0262_ ;
wire _0263_ ;
wire _0264_ ;
wire _0265_ ;
wire _0266_ ;
wire _0267_ ;
wire _0268_ ;
wire _0269_ ;
wire _0270_ ;
wire _0271_ ;
wire _0272_ ;
wire _0273_ ;
wire _0274_ ;
wire _0275_ ;
wire _0276_ ;
wire _0277_ ;
wire _0278_ ;
wire _0279_ ;
wire _0280_ ;
wire _0281_ ;
wire _0282_ ;
wire _0283_ ;
wire _0284_ ;
wire _0285_ ;
wire _0286_ ;
wire _0287_ ;
wire _0288_ ;
wire _0289_ ;
wire _0290_ ;
wire _0291_ ;
wire _0292_ ;
wire _0293_ ;
wire _0294_ ;
wire _0295_ ;
wire _0296_ ;
wire _0297_ ;
wire _0298_ ;
wire _0299_ ;
wire _0300_ ;
wire _0301_ ;
wire _0302_ ;
wire _0303_ ;
wire _0304_ ;
wire _0305_ ;
wire _0306_ ;
wire _0307_ ;
wire _0308_ ;
wire _0309_ ;
wire _0310_ ;
wire _0311_ ;
wire _0312_ ;
wire _0313_ ;
wire _0314_ ;
wire _0315_ ;
wire _0316_ ;
wire _0317_ ;
wire _0318_ ;
wire _0319_ ;
wire _0320_ ;
wire _0321_ ;
wire _0322_ ;
wire _0323_ ;
wire _0324_ ;
wire _0325_ ;
wire _0326_ ;
wire _0327_ ;
wire _0328_ ;
wire _0329_ ;
wire _0330_ ;
wire _0331_ ;
wire _0332_ ;
wire _0333_ ;
wire _0334_ ;
wire _0335_ ;
wire _0336_ ;
wire _0337_ ;
wire _0338_ ;
wire _0339_ ;
wire _0340_ ;
wire _0341_ ;
wire _0342_ ;
wire _0343_ ;
wire _0344_ ;
wire _0345_ ;
wire _0346_ ;
wire _0347_ ;
wire _0348_ ;
wire _0349_ ;
wire _0350_ ;
wire _0351_ ;
wire _0352_ ;
wire _0353_ ;
wire _0354_ ;
wire _0355_ ;
wire _0356_ ;
wire _0357_ ;
wire _0358_ ;
wire _0359_ ;
wire _0360_ ;
wire _0361_ ;
wire _0362_ ;
wire _0363_ ;
wire _0364_ ;
wire _0365_ ;
wire _0366_ ;
wire _0367_ ;
wire _0368_ ;
wire _0369_ ;
wire _0370_ ;
wire _0371_ ;
wire _0372_ ;
wire _0373_ ;
wire _0374_ ;
wire _0375_ ;
wire _0376_ ;
wire _0377_ ;
wire _0378_ ;
wire _0379_ ;
wire _0380_ ;
wire _0381_ ;
wire _0382_ ;
wire _0383_ ;
wire _0384_ ;
wire _0385_ ;
wire _0386_ ;
wire _0387_ ;
wire _0388_ ;
wire _0389_ ;
wire _0390_ ;
wire _0391_ ;
wire _0392_ ;
wire _0393_ ;
wire _0394_ ;
wire _0395_ ;
wire _0396_ ;
wire _0397_ ;
wire _0398_ ;
wire _0399_ ;
wire _0400_ ;
wire _0401_ ;
wire _0402_ ;
wire _0403_ ;
wire _0404_ ;
wire _0405_ ;
wire _0406_ ;
wire _0407_ ;
wire _0408_ ;
wire _0409_ ;
wire _0410_ ;
wire _0411_ ;
wire _0412_ ;
wire _0413_ ;
wire _0414_ ;
wire _0415_ ;
wire _0416_ ;
wire _0417_ ;
wire _0418_ ;
wire _0419_ ;
wire _0420_ ;
wire _0421_ ;
wire _0422_ ;
wire _0423_ ;
wire _0424_ ;
wire _0425_ ;
wire _0426_ ;
wire _0427_ ;
wire _0428_ ;
wire _0429_ ;
wire _0430_ ;
wire _0431_ ;
wire _0432_ ;
wire _0433_ ;
wire _0434_ ;
wire _0435_ ;
wire _0436_ ;
wire _0437_ ;
wire _0438_ ;
wire _0439_ ;
wire _0440_ ;
wire _0441_ ;
wire _0442_ ;
wire _0443_ ;
wire _0444_ ;
wire _0445_ ;
wire _0446_ ;
wire _0447_ ;
wire _0448_ ;
wire _0449_ ;
wire _0450_ ;
wire _0451_ ;
wire _0452_ ;
wire _0453_ ;
wire _0454_ ;
wire _0455_ ;
wire _0456_ ;
wire _0457_ ;
wire _0458_ ;
wire _0459_ ;
wire _0460_ ;
wire _0461_ ;
wire _0462_ ;
wire _0463_ ;
wire _0464_ ;
wire _0465_ ;
wire _0466_ ;
wire _0467_ ;
wire _0468_ ;
wire _0469_ ;
wire _0470_ ;
wire _0471_ ;
wire _0472_ ;
wire _0473_ ;
wire _0474_ ;
wire _0475_ ;
wire _0476_ ;
wire _0477_ ;
wire _0478_ ;
wire _0479_ ;
wire _0480_ ;
wire _0481_ ;
wire _0482_ ;
wire _0483_ ;
wire _0484_ ;
wire _0485_ ;
wire _0486_ ;
wire _0487_ ;
wire _0488_ ;
wire _0489_ ;
wire _0490_ ;
wire _0491_ ;
wire _0492_ ;
wire _0493_ ;
wire _0494_ ;
wire _0495_ ;
wire _0496_ ;
wire _0497_ ;
wire _0498_ ;
wire _0499_ ;
wire _0500_ ;
wire _0501_ ;
wire _0502_ ;
wire _0503_ ;
wire _0504_ ;
wire _0505_ ;
wire _0506_ ;
wire _0507_ ;
wire _0508_ ;
wire _0509_ ;
wire _0510_ ;
wire _0511_ ;
wire _0512_ ;
wire _0513_ ;
wire _0514_ ;
wire _0515_ ;
wire _0516_ ;
wire _0517_ ;
wire _0518_ ;
wire _0519_ ;
wire _0520_ ;
wire _0521_ ;
wire _0522_ ;
wire _0523_ ;
wire _0524_ ;
wire _0525_ ;
wire _0526_ ;
wire _0527_ ;
wire _0528_ ;
wire _0529_ ;
wire _0530_ ;
wire _0531_ ;
wire _0532_ ;
wire _0533_ ;
wire _0534_ ;
wire _0535_ ;
wire _0536_ ;
wire _0537_ ;
wire _0538_ ;
wire _0539_ ;
wire _0540_ ;
wire _0541_ ;
wire _0542_ ;
wire _0543_ ;
wire _0544_ ;
wire _0545_ ;
wire _0546_ ;
wire _0547_ ;
wire _0548_ ;
wire _0549_ ;
wire _0550_ ;
wire _0551_ ;
wire _0552_ ;
wire _0553_ ;
wire _0554_ ;
wire _0555_ ;
wire _0556_ ;
wire _0557_ ;
wire _0558_ ;
wire _0559_ ;
wire _0560_ ;
wire _0561_ ;
wire _0562_ ;
wire _0563_ ;
wire _0564_ ;
wire _0565_ ;
wire _0566_ ;
wire _0567_ ;
wire _0568_ ;
wire _0569_ ;
wire _0570_ ;
wire _0571_ ;
wire _0572_ ;
wire _0573_ ;
wire _0574_ ;
wire _0575_ ;
wire _0576_ ;
wire _0577_ ;
wire _0578_ ;
wire _0579_ ;
wire _0580_ ;
wire _0581_ ;
wire _0582_ ;
wire _0583_ ;
wire _0584_ ;
wire _0585_ ;
wire _0586_ ;
wire _0587_ ;
wire _0588_ ;
wire _0589_ ;
wire _0590_ ;
wire _0591_ ;
wire _0592_ ;
wire _0593_ ;
wire _0594_ ;
wire _0595_ ;
wire _0596_ ;
wire _0597_ ;
wire _0598_ ;
wire _0599_ ;
wire _0600_ ;
wire _0601_ ;
wire _0602_ ;
wire _0603_ ;
wire _0604_ ;
wire _0605_ ;
wire _0606_ ;
wire _0607_ ;
wire _0608_ ;
wire _0609_ ;
wire _0610_ ;
wire _0611_ ;
wire _0612_ ;
wire _0613_ ;
wire _0614_ ;
wire _0615_ ;
wire _0616_ ;
wire _0617_ ;
wire _0618_ ;
wire _0619_ ;
wire _0620_ ;
wire _0621_ ;
wire _0622_ ;
wire _0623_ ;
wire _0624_ ;
wire _0625_ ;
wire _0626_ ;
wire _0627_ ;
wire _0628_ ;
wire _0629_ ;
wire _0630_ ;
wire _0631_ ;
wire _0632_ ;
wire _0633_ ;
wire _0634_ ;
wire _0635_ ;
wire _0636_ ;
wire _0637_ ;
wire _0638_ ;
wire _0639_ ;
wire _0640_ ;
wire _0641_ ;
wire _0642_ ;
wire _0643_ ;
wire _0644_ ;
wire _0645_ ;
wire _0646_ ;
wire _0647_ ;
wire _0648_ ;
wire _0649_ ;
wire _0650_ ;
wire _0651_ ;
wire _0652_ ;
wire _0653_ ;
wire _0654_ ;
wire _0655_ ;
wire _0656_ ;
wire _0657_ ;
wire _0658_ ;
wire _0659_ ;
wire _0660_ ;
wire _0661_ ;
wire _0662_ ;
wire _0663_ ;
wire _0664_ ;
wire _0665_ ;
wire _0666_ ;
wire _0667_ ;
wire _0668_ ;
wire _0669_ ;
wire _0670_ ;
wire _0671_ ;
wire _0672_ ;
wire _0673_ ;
wire _0674_ ;
wire _0675_ ;
wire _0676_ ;
wire _0677_ ;
wire _0678_ ;
wire _0679_ ;
wire _0680_ ;
wire _0681_ ;
wire _0682_ ;
wire _0683_ ;
wire _0684_ ;
wire _0685_ ;
wire _0686_ ;
wire _0687_ ;
wire _0688_ ;
wire _0689_ ;
wire _0690_ ;
wire _0691_ ;
wire _0692_ ;
wire _0693_ ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XNOR__A_Y_$_NAND__A_B ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_ORNOT__Y_A_$_ORNOT__Y_B_$_XOR__A_Y_$_OR__A_1_B ;
wire ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ;
wire ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ;
wire \i0.state_$_SDFFE_PP0P__Q_E ;
wire \i0.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \inst_o[0] ;
wire \inst_o[1] ;
wire \inst_o[2] ;
wire \inst_o[3] ;
wire \inst_o[4] ;
wire \inst_o[5] ;
wire \inst_o[6] ;
wire \inst_o[7] ;
wire \inst_o[8] ;
wire \inst_o[9] ;
wire \inst_o[10] ;
wire \inst_o[11] ;
wire \inst_o[12] ;
wire \inst_o[13] ;
wire \inst_o[14] ;
wire \inst_o[15] ;
wire \inst_o[16] ;
wire \inst_o[17] ;
wire \inst_o[18] ;
wire \inst_o[19] ;
wire \inst_o[20] ;
wire \inst_o[21] ;
wire \inst_o[22] ;
wire \inst_o[23] ;
wire \inst_o[24] ;
wire \inst_o[25] ;
wire \inst_o[26] ;
wire \inst_o[27] ;
wire \inst_o[28] ;
wire \inst_o[29] ;
wire \inst_o[30] ;
wire \inst_o[31] ;
wire \i0.io_Pc_count[0] ;
wire \i0.io_Pc_count[1] ;
wire \i0.io_Pc_count[2] ;
wire \i0.io_Pc_count[3] ;
wire \i0.io_Pc_count[4] ;
wire \i0.io_Pc_count[5] ;
wire \i0.io_Pc_count[6] ;
wire \i0.io_Pc_count[7] ;
wire \i0.io_Pc_count[8] ;
wire \i0.io_Pc_count[9] ;
wire \i0.io_Pc_count[10] ;
wire \i0.io_Pc_count[11] ;
wire \i0.io_Pc_count[12] ;
wire \i0.io_Pc_count[13] ;
wire \i0.io_Pc_count[14] ;
wire \i0.io_Pc_count[15] ;
wire \i0.io_Pc_count[16] ;
wire \i0.io_Pc_count[17] ;
wire \i0.io_Pc_count[18] ;
wire \i0.io_Pc_count[19] ;
wire \i0.io_Pc_count[20] ;
wire \i0.io_Pc_count[21] ;
wire \i0.io_Pc_count[22] ;
wire \i0.io_Pc_count[23] ;
wire \i0.io_Pc_count[24] ;
wire \i0.io_Pc_count[25] ;
wire \i0.io_Pc_count[26] ;
wire \i0.io_Pc_count[27] ;
wire \i0.io_Pc_count[28] ;
wire \i0.io_Pc_count[29] ;
wire \i0.io_Pc_count[30] ;
wire \i0.io_Pc_count[31] ;
wire \i5.io_mem_data[0] ;
wire \i5.io_mem_data[1] ;
wire \i5.io_mem_data[2] ;
wire \i5.io_mem_data[3] ;
wire \i5.io_mem_data[4] ;
wire \i5.io_mem_data[5] ;
wire \i5.io_mem_data[6] ;
wire \i5.io_mem_data[7] ;

assign inst_o[0] = \inst_o[0] ;
assign inst_o[0] = \inst_o[1] ;
assign inst_o[2] = \inst_o[2] ;
assign inst_o[3] = \inst_o[3] ;
assign inst_o[4] = \inst_o[4] ;
assign inst_o[5] = \inst_o[5] ;
assign inst_o[6] = \inst_o[6] ;
assign inst_o[7] = \inst_o[7] ;
assign inst_o[10] = \inst_o[8] ;
assign inst_o[10] = \inst_o[9] ;
assign inst_o[10] = \inst_o[10] ;
assign inst_o[10] = \inst_o[11] ;
assign inst_o[10] = \inst_o[12] ;
assign inst_o[10] = \inst_o[13] ;
assign inst_o[10] = \inst_o[14] ;
assign inst_o[10] = \inst_o[15] ;
assign inst_o[10] = \inst_o[16] ;
assign inst_o[10] = \inst_o[17] ;
assign inst_o[10] = \inst_o[18] ;
assign inst_o[10] = \inst_o[19] ;
assign inst_o[10] = \inst_o[20] ;
assign inst_o[10] = \inst_o[21] ;
assign inst_o[10] = \inst_o[22] ;
assign inst_o[10] = \inst_o[23] ;
assign inst_o[10] = \inst_o[24] ;
assign inst_o[10] = \inst_o[25] ;
assign inst_o[10] = \inst_o[26] ;
assign inst_o[10] = \inst_o[27] ;
assign inst_o[10] = \inst_o[28] ;
assign inst_o[10] = \inst_o[29] ;
assign inst_o[10] = \inst_o[30] ;
assign inst_o[10] = \inst_o[31] ;

INV_X32 _0694_ ( .A(\inst_o[5] ), .ZN(_0044_ ) );
NOR2_X4 _0695_ ( .A1(_0044_ ), .A2(\inst_o[4] ), .ZN(_0045_ ) );
AND2_X4 _0696_ ( .A1(_0045_ ), .A2(\inst_o[6] ), .ZN(_0046_ ) );
INV_X1 _0697_ ( .A(_0046_ ), .ZN(_0047_ ) );
INV_X1 _0698_ ( .A(\inst_o[3] ), .ZN(_0048_ ) );
NAND3_X1 _0699_ ( .A1(_0048_ ), .A2(\inst_o[2] ), .A3(\inst_o[0] ), .ZN(_0049_ ) );
NOR2_X1 _0700_ ( .A1(_0047_ ), .A2(_0049_ ), .ZN(_0050_ ) );
NOR2_X1 _0701_ ( .A1(_0050_ ), .A2(reset ), .ZN(_0051_ ) );
NOR2_X1 _0702_ ( .A1(\inst_o[3] ), .A2(\inst_o[2] ), .ZN(_0052_ ) );
AND2_X2 _0703_ ( .A1(_0052_ ), .A2(\inst_o[0] ), .ZN(_0053_ ) );
AND2_X1 _0704_ ( .A1(_0046_ ), .A2(_0053_ ), .ZN(_0054_ ) );
INV_X1 _0705_ ( .A(_0054_ ), .ZN(_0055_ ) );
BUF_X2 _0706_ ( .A(_0055_ ), .Z(_0056_ ) );
INV_X1 _0707_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0057_ ) );
AND2_X2 _0708_ ( .A1(\i0.io_Pc_count[3] ), .A2(\i0.io_Pc_count[2] ), .ZN(_0058_ ) );
AND2_X1 _0709_ ( .A1(\i0.io_Pc_count[5] ), .A2(\i0.io_Pc_count[4] ), .ZN(_0059_ ) );
AND2_X1 _0710_ ( .A1(\i0.io_Pc_count[7] ), .A2(\i0.io_Pc_count[6] ), .ZN(_0060_ ) );
AND4_X1 _0711_ ( .A1(\i0.io_Pc_count[9] ), .A2(_0058_ ), .A3(_0059_ ), .A4(_0060_ ), .ZN(_0061_ ) );
AND2_X1 _0712_ ( .A1(_0061_ ), .A2(\i0.io_Pc_count[8] ), .ZN(_0062_ ) );
OAI211_X1 _0713_ ( .A(_0051_ ), .B(_0056_ ), .C1(_0057_ ), .C2(_0062_ ), .ZN(_0063_ ) );
AND2_X1 _0714_ ( .A1(_0062_ ), .A2(_0057_ ), .ZN(_0064_ ) );
NOR2_X1 _0715_ ( .A1(_0063_ ), .A2(_0064_ ), .ZN(_0000_ ) );
AND2_X1 _0716_ ( .A1(_0058_ ), .A2(_0059_ ), .ZN(_0065_ ) );
AND2_X1 _0717_ ( .A1(_0065_ ), .A2(_0060_ ), .ZN(_0066_ ) );
INV_X1 _0718_ ( .A(_0066_ ), .ZN(_0067_ ) );
NOR2_X1 _0719_ ( .A1(_0067_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0068_ ) );
XOR2_X1 _0720_ ( .A(_0068_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .Z(_0069_ ) );
NAND2_X1 _0721_ ( .A1(_0051_ ), .A2(_0056_ ), .ZN(_0070_ ) );
NOR2_X1 _0722_ ( .A1(_0069_ ), .A2(_0070_ ), .ZN(_0001_ ) );
INV_X1 _0723_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0071_ ) );
NAND4_X1 _0724_ ( .A1(_0071_ ), .A2(\inst_o[7] ), .A3(\i0.io_Pc_count[14] ), .A4(\i0.io_Pc_count[11] ), .ZN(_0072_ ) );
INV_X1 _0725_ ( .A(\i0.io_Pc_count[13] ), .ZN(_0073_ ) );
NOR2_X1 _0726_ ( .A1(_0072_ ), .A2(_0073_ ), .ZN(_0074_ ) );
AND2_X1 _0727_ ( .A1(\i0.io_Pc_count[15] ), .A2(\i0.io_Pc_count[16] ), .ZN(_0075_ ) );
AND2_X2 _0728_ ( .A1(_0074_ ), .A2(_0075_ ), .ZN(_0076_ ) );
AND3_X1 _0729_ ( .A1(\i0.io_Pc_count[19] ), .A2(\i0.io_Pc_count[18] ), .A3(\i0.io_Pc_count[17] ), .ZN(_0077_ ) );
AND2_X2 _0730_ ( .A1(_0077_ ), .A2(\i0.io_Pc_count[20] ), .ZN(_0078_ ) );
AND3_X1 _0731_ ( .A1(\i0.io_Pc_count[23] ), .A2(\i0.io_Pc_count[22] ), .A3(\i0.io_Pc_count[21] ), .ZN(_0079_ ) );
AND2_X1 _0732_ ( .A1(_0079_ ), .A2(\i0.io_Pc_count[24] ), .ZN(_0080_ ) );
AND2_X1 _0733_ ( .A1(\i0.io_Pc_count[26] ), .A2(\i0.io_Pc_count[25] ), .ZN(_0081_ ) );
AND3_X1 _0734_ ( .A1(_0081_ ), .A2(\i0.io_Pc_count[28] ), .A3(\i0.io_Pc_count[27] ), .ZN(_0082_ ) );
NAND4_X1 _0735_ ( .A1(_0076_ ), .A2(_0078_ ), .A3(_0080_ ), .A4(_0082_ ), .ZN(_0083_ ) );
BUF_X4 _0736_ ( .A(_0054_ ), .Z(_0084_ ) );
MUX2_X1 _0737_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .B(_0083_ ), .S(_0084_ ), .Z(_0085_ ) );
AND3_X1 _0738_ ( .A1(_0062_ ), .A2(\i0.io_Pc_count[11] ), .A3(\i0.io_Pc_count[10] ), .ZN(_0086_ ) );
AND4_X1 _0739_ ( .A1(\i0.io_Pc_count[15] ), .A2(_0086_ ), .A3(\i0.io_Pc_count[13] ), .A4(\i0.io_Pc_count[12] ), .ZN(_0087_ ) );
AND3_X1 _0740_ ( .A1(_0087_ ), .A2(\i0.io_Pc_count[16] ), .A3(\i0.io_Pc_count[14] ), .ZN(_0088_ ) );
AND3_X1 _0741_ ( .A1(_0088_ ), .A2(\i0.io_Pc_count[20] ), .A3(_0077_ ), .ZN(_0089_ ) );
AND3_X1 _0742_ ( .A1(\i0.io_Pc_count[27] ), .A2(\i0.io_Pc_count[26] ), .A3(\i0.io_Pc_count[25] ), .ZN(_0090_ ) );
NAND4_X1 _0743_ ( .A1(_0089_ ), .A2(\i0.io_Pc_count[24] ), .A3(_0090_ ), .A4(_0079_ ), .ZN(_0091_ ) );
AOI21_X1 _0744_ ( .A(_0085_ ), .B1(_0091_ ), .B2(_0056_ ), .ZN(_0092_ ) );
XNOR2_X1 _0745_ ( .A(_0092_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0093_ ) );
AND2_X1 _0746_ ( .A1(_0093_ ), .A2(_0051_ ), .ZN(_0002_ ) );
AND2_X1 _0747_ ( .A1(\i0.io_Pc_count[11] ), .A2(\i0.io_Pc_count[10] ), .ZN(_0094_ ) );
AND2_X1 _0748_ ( .A1(_0062_ ), .A2(_0094_ ), .ZN(_0095_ ) );
AND3_X1 _0749_ ( .A1(_0095_ ), .A2(\i0.io_Pc_count[13] ), .A3(\i0.io_Pc_count[12] ), .ZN(_0096_ ) );
AND3_X1 _0750_ ( .A1(_0096_ ), .A2(\i0.io_Pc_count[15] ), .A3(\i0.io_Pc_count[14] ), .ZN(_0097_ ) );
AND3_X1 _0751_ ( .A1(_0097_ ), .A2(\i0.io_Pc_count[16] ), .A3(_0078_ ), .ZN(_0098_ ) );
BUF_X2 _0752_ ( .A(_0080_ ), .Z(_0099_ ) );
NAND4_X1 _0753_ ( .A1(_0098_ ), .A2(_0056_ ), .A3(_0090_ ), .A4(_0099_ ), .ZN(_0100_ ) );
AND2_X1 _0754_ ( .A1(_0054_ ), .A2(_0076_ ), .ZN(_0101_ ) );
AND2_X1 _0755_ ( .A1(_0101_ ), .A2(_0078_ ), .ZN(_0102_ ) );
INV_X1 _0756_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0103_ ) );
NAND4_X1 _0757_ ( .A1(_0102_ ), .A2(_0103_ ), .A3(_0081_ ), .A4(_0099_ ), .ZN(_0104_ ) );
AND3_X1 _0758_ ( .A1(_0100_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_0104_ ), .ZN(_0105_ ) );
AOI21_X1 _0759_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0100_ ), .B2(_0104_ ), .ZN(_0106_ ) );
INV_X1 _0760_ ( .A(_0051_ ), .ZN(_0107_ ) );
BUF_X4 _0761_ ( .A(_0107_ ), .Z(_0108_ ) );
NOR3_X1 _0762_ ( .A1(_0105_ ), .A2(_0106_ ), .A3(_0108_ ), .ZN(_0003_ ) );
NAND3_X1 _0763_ ( .A1(_0098_ ), .A2(\i0.io_Pc_count[25] ), .A3(_0099_ ), .ZN(_0109_ ) );
AND2_X1 _0764_ ( .A1(_0109_ ), .A2(_0056_ ), .ZN(_0110_ ) );
NAND3_X1 _0765_ ( .A1(_0102_ ), .A2(_0081_ ), .A3(_0099_ ), .ZN(_0111_ ) );
INV_X1 _0766_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0112_ ) );
INV_X1 _0767_ ( .A(_0053_ ), .ZN(_0113_ ) );
OAI21_X1 _0768_ ( .A(_0112_ ), .B1(_0047_ ), .B2(_0113_ ), .ZN(_0114_ ) );
AOI21_X1 _0769_ ( .A(_0110_ ), .B1(_0111_ ), .B2(_0114_ ), .ZN(_0115_ ) );
AND2_X1 _0770_ ( .A1(_0115_ ), .A2(_0103_ ), .ZN(_0116_ ) );
NOR2_X1 _0771_ ( .A1(_0115_ ), .A2(_0103_ ), .ZN(_0117_ ) );
NOR3_X1 _0772_ ( .A1(_0116_ ), .A2(_0117_ ), .A3(_0108_ ), .ZN(_0004_ ) );
NAND4_X1 _0773_ ( .A1(_0098_ ), .A2(\i0.io_Pc_count[25] ), .A3(_0056_ ), .A4(_0099_ ), .ZN(_0118_ ) );
NAND2_X1 _0774_ ( .A1(_0102_ ), .A2(_0099_ ), .ZN(_0119_ ) );
OR2_X1 _0775_ ( .A1(_0119_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0120_ ) );
NAND2_X1 _0776_ ( .A1(_0118_ ), .A2(_0120_ ), .ZN(_0121_ ) );
OAI21_X1 _0777_ ( .A(_0051_ ), .B1(_0121_ ), .B2(_0112_ ), .ZN(_0122_ ) );
AOI21_X1 _0778_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0118_ ), .B2(_0120_ ), .ZN(_0123_ ) );
NOR2_X1 _0779_ ( .A1(_0122_ ), .A2(_0123_ ), .ZN(_0005_ ) );
NAND4_X1 _0780_ ( .A1(_0084_ ), .A2(_0076_ ), .A3(_0078_ ), .A4(_0099_ ), .ZN(_0124_ ) );
BUF_X4 _0781_ ( .A(_0084_ ), .Z(_0125_ ) );
OAI21_X1 _0782_ ( .A(_0124_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .B2(_0125_ ), .ZN(_0126_ ) );
AND2_X1 _0783_ ( .A1(_0098_ ), .A2(_0079_ ), .ZN(_0127_ ) );
OAI21_X1 _0784_ ( .A(_0126_ ), .B1(_0127_ ), .B2(_0125_ ), .ZN(_0128_ ) );
AND2_X1 _0785_ ( .A1(_0128_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0129_ ) );
NOR2_X1 _0786_ ( .A1(_0128_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0130_ ) );
NOR3_X1 _0787_ ( .A1(_0129_ ), .A2(_0130_ ), .A3(_0108_ ), .ZN(_0006_ ) );
AND2_X1 _0788_ ( .A1(_0097_ ), .A2(\i0.io_Pc_count[16] ), .ZN(_0131_ ) );
NAND4_X1 _0789_ ( .A1(_0131_ ), .A2(_0055_ ), .A3(_0078_ ), .A4(_0079_ ), .ZN(_0132_ ) );
INV_X1 _0790_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0133_ ) );
AND2_X1 _0791_ ( .A1(\i0.io_Pc_count[22] ), .A2(\i0.io_Pc_count[21] ), .ZN(_0134_ ) );
NAND4_X1 _0792_ ( .A1(_0101_ ), .A2(_0133_ ), .A3(_0078_ ), .A4(_0134_ ), .ZN(_0135_ ) );
AND2_X1 _0793_ ( .A1(_0132_ ), .A2(_0135_ ), .ZN(_0136_ ) );
OR2_X1 _0794_ ( .A1(_0136_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0137_ ) );
AOI21_X1 _0795_ ( .A(_0107_ ), .B1(_0136_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0138_ ) );
AND2_X1 _0796_ ( .A1(_0137_ ), .A2(_0138_ ), .ZN(_0007_ ) );
AOI21_X1 _0797_ ( .A(_0084_ ), .B1(_0098_ ), .B2(\i0.io_Pc_count[21] ), .ZN(_0139_ ) );
NAND3_X1 _0798_ ( .A1(_0101_ ), .A2(_0078_ ), .A3(_0134_ ), .ZN(_0140_ ) );
INV_X1 _0799_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0141_ ) );
OAI21_X1 _0800_ ( .A(_0141_ ), .B1(_0047_ ), .B2(_0113_ ), .ZN(_0142_ ) );
AOI21_X1 _0801_ ( .A(_0139_ ), .B1(_0140_ ), .B2(_0142_ ), .ZN(_0143_ ) );
AND2_X1 _0802_ ( .A1(_0143_ ), .A2(_0133_ ), .ZN(_0144_ ) );
NOR2_X1 _0803_ ( .A1(_0143_ ), .A2(_0133_ ), .ZN(_0145_ ) );
NOR3_X1 _0804_ ( .A1(_0144_ ), .A2(_0145_ ), .A3(_0108_ ), .ZN(_0008_ ) );
NAND4_X1 _0805_ ( .A1(_0131_ ), .A2(\i0.io_Pc_count[21] ), .A3(_0056_ ), .A4(_0078_ ), .ZN(_0146_ ) );
INV_X1 _0806_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0147_ ) );
NAND4_X1 _0807_ ( .A1(_0125_ ), .A2(_0076_ ), .A3(_0147_ ), .A4(_0078_ ), .ZN(_0148_ ) );
NAND2_X1 _0808_ ( .A1(_0146_ ), .A2(_0148_ ), .ZN(_0149_ ) );
OAI21_X1 _0809_ ( .A(_0051_ ), .B1(_0149_ ), .B2(_0141_ ), .ZN(_0150_ ) );
AOI21_X1 _0810_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0146_ ), .B2(_0148_ ), .ZN(_0151_ ) );
NOR2_X1 _0811_ ( .A1(_0150_ ), .A2(_0151_ ), .ZN(_0009_ ) );
AOI21_X1 _0812_ ( .A(_0084_ ), .B1(_0088_ ), .B2(_0077_ ), .ZN(_0152_ ) );
INV_X1 _0813_ ( .A(_0102_ ), .ZN(_0153_ ) );
OR2_X1 _0814_ ( .A1(_0084_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0154_ ) );
AOI21_X1 _0815_ ( .A(_0152_ ), .B1(_0153_ ), .B2(_0154_ ), .ZN(_0155_ ) );
AND2_X1 _0816_ ( .A1(_0155_ ), .A2(_0147_ ), .ZN(_0156_ ) );
NOR2_X1 _0817_ ( .A1(_0155_ ), .A2(_0147_ ), .ZN(_0157_ ) );
NOR3_X1 _0818_ ( .A1(_0156_ ), .A2(_0157_ ), .A3(_0108_ ), .ZN(_0010_ ) );
NAND4_X1 _0819_ ( .A1(_0097_ ), .A2(\i0.io_Pc_count[16] ), .A3(_0055_ ), .A4(_0077_ ), .ZN(_0158_ ) );
NAND3_X1 _0820_ ( .A1(_0101_ ), .A2(\i0.io_Pc_count[18] ), .A3(\i0.io_Pc_count[17] ), .ZN(_0159_ ) );
OR2_X1 _0821_ ( .A1(_0159_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0160_ ) );
AND2_X1 _0822_ ( .A1(_0158_ ), .A2(_0160_ ), .ZN(_0161_ ) );
OR2_X1 _0823_ ( .A1(_0161_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0162_ ) );
AOI21_X1 _0824_ ( .A(_0107_ ), .B1(_0161_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0163_ ) );
AND2_X1 _0825_ ( .A1(_0162_ ), .A2(_0163_ ), .ZN(_0011_ ) );
AOI21_X1 _0826_ ( .A(_0070_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .B2(_0067_ ), .ZN(_0164_ ) );
INV_X1 _0827_ ( .A(_0068_ ), .ZN(_0165_ ) );
AND2_X1 _0828_ ( .A1(_0164_ ), .A2(_0165_ ), .ZN(_0012_ ) );
NAND4_X1 _0829_ ( .A1(_0084_ ), .A2(_0076_ ), .A3(\i0.io_Pc_count[18] ), .A4(\i0.io_Pc_count[17] ), .ZN(_0166_ ) );
OAI21_X1 _0830_ ( .A(_0166_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .B2(_0084_ ), .ZN(_0167_ ) );
AND4_X1 _0831_ ( .A1(\i0.io_Pc_count[16] ), .A2(_0087_ ), .A3(\i0.io_Pc_count[17] ), .A4(\i0.io_Pc_count[14] ), .ZN(_0168_ ) );
OAI21_X1 _0832_ ( .A(_0167_ ), .B1(_0168_ ), .B2(_0125_ ), .ZN(_0169_ ) );
AND2_X1 _0833_ ( .A1(_0169_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0170_ ) );
NOR2_X1 _0834_ ( .A1(_0169_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0171_ ) );
NOR3_X1 _0835_ ( .A1(_0170_ ), .A2(_0171_ ), .A3(_0108_ ), .ZN(_0013_ ) );
NAND4_X1 _0836_ ( .A1(_0097_ ), .A2(\i0.io_Pc_count[16] ), .A3(\i0.io_Pc_count[17] ), .A4(_0056_ ), .ZN(_0172_ ) );
INV_X1 _0837_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0173_ ) );
NAND3_X1 _0838_ ( .A1(_0125_ ), .A2(_0076_ ), .A3(_0173_ ), .ZN(_0174_ ) );
AND3_X1 _0839_ ( .A1(_0172_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_0174_ ), .ZN(_0175_ ) );
AOI21_X1 _0840_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0172_ ), .B2(_0174_ ), .ZN(_0176_ ) );
NOR3_X1 _0841_ ( .A1(_0175_ ), .A2(_0176_ ), .A3(_0108_ ), .ZN(_0014_ ) );
AOI21_X1 _0842_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0046_ ), .B2(_0053_ ), .ZN(_0177_ ) );
NAND4_X1 _0843_ ( .A1(_0096_ ), .A2(\i0.io_Pc_count[15] ), .A3(\i0.io_Pc_count[14] ), .A4(_0177_ ), .ZN(_0178_ ) );
INV_X1 _0844_ ( .A(_0101_ ), .ZN(_0179_ ) );
AND3_X1 _0845_ ( .A1(_0178_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_0179_ ), .ZN(_0180_ ) );
AOI21_X1 _0846_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0178_ ), .B2(_0179_ ), .ZN(_0181_ ) );
NOR3_X1 _0847_ ( .A1(_0180_ ), .A2(_0181_ ), .A3(_0108_ ), .ZN(_0015_ ) );
NAND4_X1 _0848_ ( .A1(_0096_ ), .A2(\i0.io_Pc_count[15] ), .A3(\i0.io_Pc_count[14] ), .A4(_0055_ ), .ZN(_0182_ ) );
INV_X1 _0849_ ( .A(_0074_ ), .ZN(_0183_ ) );
OR4_X1 _0850_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(_0047_ ), .A3(_0183_ ), .A4(_0113_ ), .ZN(_0184_ ) );
AND2_X1 _0851_ ( .A1(_0182_ ), .A2(_0184_ ), .ZN(_0185_ ) );
OR2_X1 _0852_ ( .A1(_0185_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0186_ ) );
AOI21_X1 _0853_ ( .A(_0107_ ), .B1(_0185_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0187_ ) );
AND2_X1 _0854_ ( .A1(_0186_ ), .A2(_0187_ ), .ZN(_0016_ ) );
OR2_X1 _0855_ ( .A1(_0096_ ), .A2(_0084_ ), .ZN(_0188_ ) );
AND3_X1 _0856_ ( .A1(_0046_ ), .A2(_0074_ ), .A3(_0053_ ), .ZN(_0189_ ) );
AOI21_X1 _0857_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_0046_ ), .B2(_0053_ ), .ZN(_0190_ ) );
OAI21_X1 _0858_ ( .A(_0188_ ), .B1(_0189_ ), .B2(_0190_ ), .ZN(_0191_ ) );
AND2_X1 _0859_ ( .A1(_0191_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0192_ ) );
NOR2_X1 _0860_ ( .A1(_0191_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0193_ ) );
NOR3_X1 _0861_ ( .A1(_0192_ ), .A2(_0193_ ), .A3(_0108_ ), .ZN(_0017_ ) );
AND2_X1 _0862_ ( .A1(\inst_o[7] ), .A2(\i0.io_Pc_count[11] ), .ZN(_0194_ ) );
AND2_X1 _0863_ ( .A1(_0194_ ), .A2(_0071_ ), .ZN(_0195_ ) );
OR3_X1 _0864_ ( .A1(_0047_ ), .A2(_0113_ ), .A3(_0195_ ), .ZN(_0196_ ) );
NAND4_X1 _0865_ ( .A1(_0053_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\inst_o[6] ), .A4(_0045_ ), .ZN(_0197_ ) );
NAND3_X1 _0866_ ( .A1(_0188_ ), .A2(_0196_ ), .A3(_0197_ ), .ZN(_0198_ ) );
OAI21_X1 _0867_ ( .A(_0051_ ), .B1(_0198_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0199_ ) );
AOI21_X1 _0868_ ( .A(_0199_ ), .B1(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .B2(_0198_ ), .ZN(_0018_ ) );
MUX2_X1 _0869_ ( .A(_0194_ ), .B(_0095_ ), .S(_0055_ ), .Z(_0200_ ) );
INV_X1 _0870_ ( .A(_0200_ ), .ZN(_0201_ ) );
OR2_X1 _0871_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0202_ ) );
NOR2_X1 _0872_ ( .A1(_0201_ ), .A2(_0202_ ), .ZN(_0203_ ) );
AND2_X1 _0873_ ( .A1(_0200_ ), .A2(_0071_ ), .ZN(_0204_ ) );
INV_X1 _0874_ ( .A(_0204_ ), .ZN(_0205_ ) );
AOI211_X1 _0875_ ( .A(_0108_ ), .B(_0203_ ), .C1(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .C2(_0205_ ), .ZN(_0019_ ) );
OAI21_X1 _0876_ ( .A(_0051_ ), .B1(_0200_ ), .B2(_0071_ ), .ZN(_0206_ ) );
NOR2_X1 _0877_ ( .A1(_0204_ ), .A2(_0206_ ), .ZN(_0020_ ) );
XNOR2_X1 _0878_ ( .A(\inst_o[7] ), .B(\i0.io_Pc_count[11] ), .ZN(_0207_ ) );
AND4_X1 _0879_ ( .A1(\inst_o[6] ), .A2(_0053_ ), .A3(_0045_ ), .A4(_0207_ ), .ZN(_0208_ ) );
XOR2_X1 _0880_ ( .A(_0064_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .Z(_0209_ ) );
AOI211_X1 _0881_ ( .A(_0107_ ), .B(_0208_ ), .C1(_0209_ ), .C2(_0056_ ), .ZN(_0021_ ) );
INV_X1 _0882_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0210_ ) );
NAND3_X1 _0883_ ( .A1(_0058_ ), .A2(_0059_ ), .A3(_0210_ ), .ZN(_0211_ ) );
XNOR2_X1 _0884_ ( .A(_0211_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0212_ ) );
NOR4_X1 _0885_ ( .A1(_0212_ ), .A2(_0050_ ), .A3(_0125_ ), .A4(reset ), .ZN(_0022_ ) );
XNOR2_X1 _0886_ ( .A(_0065_ ), .B(_0210_ ), .ZN(_0213_ ) );
NOR4_X1 _0887_ ( .A1(_0213_ ), .A2(_0050_ ), .A3(_0125_ ), .A4(reset ), .ZN(_0023_ ) );
INV_X1 _0888_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0214_ ) );
INV_X1 _0889_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0215_ ) );
AOI21_X1 _0890_ ( .A(_0214_ ), .B1(_0058_ ), .B2(_0215_ ), .ZN(_0216_ ) );
AND4_X1 _0891_ ( .A1(\i0.io_Pc_count[3] ), .A2(_0214_ ), .A3(_0215_ ), .A4(\i0.io_Pc_count[2] ), .ZN(_0217_ ) );
NOR3_X1 _0892_ ( .A1(_0070_ ), .A2(_0216_ ), .A3(_0217_ ), .ZN(_0024_ ) );
XNOR2_X1 _0893_ ( .A(_0058_ ), .B(_0215_ ), .ZN(_0218_ ) );
NOR4_X1 _0894_ ( .A1(_0050_ ), .A2(_0125_ ), .A3(reset ), .A4(_0218_ ), .ZN(_0025_ ) );
NOR2_X1 _0895_ ( .A1(\i0.io_Pc_count[3] ), .A2(\i0.io_Pc_count[2] ), .ZN(_0219_ ) );
NOR3_X1 _0896_ ( .A1(_0070_ ), .A2(_0058_ ), .A3(_0219_ ), .ZN(_0026_ ) );
NOR4_X1 _0897_ ( .A1(_0050_ ), .A2(_0125_ ), .A3(reset ), .A4(\i0.io_Pc_count[2] ), .ZN(_0027_ ) );
AND2_X1 _0898_ ( .A1(_0098_ ), .A2(_0099_ ), .ZN(_0220_ ) );
AND2_X1 _0899_ ( .A1(_0082_ ), .A2(\i0.io_Pc_count[29] ), .ZN(_0221_ ) );
NAND3_X1 _0900_ ( .A1(_0220_ ), .A2(_0056_ ), .A3(_0221_ ), .ZN(_0222_ ) );
NAND3_X1 _0901_ ( .A1(_0102_ ), .A2(_0099_ ), .A3(_0082_ ), .ZN(_0223_ ) );
OR2_X1 _0902_ ( .A1(_0223_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0224_ ) );
NAND2_X1 _0903_ ( .A1(_0222_ ), .A2(_0224_ ), .ZN(_0225_ ) );
INV_X1 _0904_ ( .A(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_0226_ ) );
OAI21_X1 _0905_ ( .A(_0051_ ), .B1(_0225_ ), .B2(_0226_ ), .ZN(_0227_ ) );
AOI21_X1 _0906_ ( .A(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .B1(_0222_ ), .B2(_0224_ ), .ZN(_0228_ ) );
NOR2_X1 _0907_ ( .A1(_0227_ ), .A2(_0228_ ), .ZN(_0028_ ) );
NAND4_X1 _0908_ ( .A1(_0220_ ), .A2(_0226_ ), .A3(_0055_ ), .A4(_0221_ ), .ZN(_0229_ ) );
AND4_X1 _0909_ ( .A1(\i0.io_Pc_count[30] ), .A2(_0084_ ), .A3(_0078_ ), .A4(_0099_ ), .ZN(_0230_ ) );
AND4_X1 _0910_ ( .A1(\i0.io_Pc_count[29] ), .A2(_0074_ ), .A3(_0082_ ), .A4(_0075_ ), .ZN(_0231_ ) );
NAND2_X1 _0911_ ( .A1(_0230_ ), .A2(_0231_ ), .ZN(_0232_ ) );
AND3_X1 _0912_ ( .A1(_0229_ ), .A2(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(_0232_ ), .ZN(_0233_ ) );
AOI21_X1 _0913_ ( .A(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_0229_ ), .B2(_0232_ ), .ZN(_0234_ ) );
NOR4_X1 _0914_ ( .A1(_0233_ ), .A2(_0234_ ), .A3(reset ), .A4(_0050_ ), .ZN(_0235_ ) );
OR2_X1 _0915_ ( .A1(_0235_ ), .A2(reset ), .ZN(_0029_ ) );
INV_X1 _0916_ ( .A(\i0.io_Pc_count[7] ), .ZN(_0236_ ) );
NOR2_X1 _0917_ ( .A1(_0236_ ), .A2(reset ), .ZN(_0030_ ) );
INV_X1 _0918_ ( .A(\i0.io_Pc_count[6] ), .ZN(_0237_ ) );
NOR2_X1 _0919_ ( .A1(_0237_ ), .A2(reset ), .ZN(_0031_ ) );
INV_X1 _0920_ ( .A(\i0.io_Pc_count[5] ), .ZN(_0238_ ) );
NOR2_X1 _0921_ ( .A1(_0238_ ), .A2(reset ), .ZN(_0032_ ) );
INV_X1 _0922_ ( .A(\i0.io_Pc_count[4] ), .ZN(_0239_ ) );
NOR2_X1 _0923_ ( .A1(_0239_ ), .A2(reset ), .ZN(_0033_ ) );
INV_X1 _0924_ ( .A(\i0.io_Pc_count[3] ), .ZN(_0240_ ) );
NOR2_X1 _0925_ ( .A1(_0240_ ), .A2(reset ), .ZN(_0034_ ) );
INV_X1 _0926_ ( .A(\i0.io_Pc_count[2] ), .ZN(_0241_ ) );
NOR2_X1 _0927_ ( .A1(_0241_ ), .A2(reset ), .ZN(_0035_ ) );
AND2_X1 _0928_ ( .A1(\inst_o[2] ), .A2(\inst_o[0] ), .ZN(_0242_ ) );
AND2_X4 _0929_ ( .A1(_0046_ ), .A2(_0242_ ), .ZN(_0243_ ) );
INV_X1 _0930_ ( .A(\inst_o[2] ), .ZN(_0244_ ) );
NOR2_X4 _0931_ ( .A1(_0243_ ), .A2(_0244_ ), .ZN(_0245_ ) );
INV_X1 _0932_ ( .A(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XNOR__A_Y_$_NAND__A_B ), .ZN(_0246_ ) );
NOR2_X1 _0933_ ( .A1(_0245_ ), .A2(_0246_ ), .ZN(_0247_ ) );
BUF_X2 _0934_ ( .A(_0247_ ), .Z(_0248_ ) );
INV_X1 _0935_ ( .A(\inst_o[0] ), .ZN(_0249_ ) );
AND2_X2 _0936_ ( .A1(_0248_ ), .A2(_0249_ ), .ZN(_0250_ ) );
AND2_X1 _0937_ ( .A1(\inst_o[6] ), .A2(\inst_o[7] ), .ZN(_0251_ ) );
AND2_X1 _0938_ ( .A1(\inst_o[4] ), .A2(\inst_o[5] ), .ZN(_0252_ ) );
AND2_X1 _0939_ ( .A1(_0251_ ), .A2(_0252_ ), .ZN(_0253_ ) );
NAND2_X1 _0940_ ( .A1(_0250_ ), .A2(_0253_ ), .ZN(_0254_ ) );
AND2_X4 _0941_ ( .A1(_0245_ ), .A2(_0246_ ), .ZN(_0255_ ) );
AND2_X1 _0942_ ( .A1(_0255_ ), .A2(_0249_ ), .ZN(_0256_ ) );
CLKBUF_X2 _0943_ ( .A(_0256_ ), .Z(_0257_ ) );
INV_X1 _0944_ ( .A(_0257_ ), .ZN(_0258_ ) );
AND2_X2 _0945_ ( .A1(_0045_ ), .A2(_0251_ ), .ZN(_0259_ ) );
INV_X1 _0946_ ( .A(_0259_ ), .ZN(_0260_ ) );
OAI21_X1 _0947_ ( .A(_0254_ ), .B1(_0258_ ), .B2(_0260_ ), .ZN(_0261_ ) );
AND2_X1 _0948_ ( .A1(_0257_ ), .A2(_0253_ ), .ZN(_0262_ ) );
NOR2_X4 _0949_ ( .A1(_0245_ ), .A2(_0048_ ), .ZN(_0263_ ) );
INV_X1 _0950_ ( .A(\inst_o[7] ), .ZN(_0264_ ) );
NOR2_X4 _0951_ ( .A1(_0264_ ), .A2(\inst_o[6] ), .ZN(_0265_ ) );
NAND4_X1 _0952_ ( .A1(_0045_ ), .A2(_0265_ ), .A3(\inst_o[0] ), .A4(_0052_ ), .ZN(_0266_ ) );
AND2_X1 _0953_ ( .A1(_0266_ ), .A2(\inst_o[0] ), .ZN(_0267_ ) );
INV_X1 _0954_ ( .A(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_ORNOT__Y_A_$_ORNOT__Y_B_$_XOR__A_Y_$_OR__A_1_B ), .ZN(_0268_ ) );
AND2_X4 _0955_ ( .A1(_0267_ ), .A2(_0268_ ), .ZN(_0269_ ) );
AND2_X1 _0956_ ( .A1(_0263_ ), .A2(_0269_ ), .ZN(_0270_ ) );
AND2_X1 _0957_ ( .A1(_0270_ ), .A2(_0253_ ), .ZN(_0271_ ) );
NOR3_X1 _0958_ ( .A1(_0261_ ), .A2(_0262_ ), .A3(_0271_ ), .ZN(_0272_ ) );
AND2_X4 _0959_ ( .A1(_0255_ ), .A2(_0269_ ), .ZN(_0273_ ) );
INV_X1 _0960_ ( .A(_0273_ ), .ZN(_0274_ ) );
AND2_X1 _0961_ ( .A1(_0044_ ), .A2(\inst_o[4] ), .ZN(_0275_ ) );
AND2_X1 _0962_ ( .A1(_0275_ ), .A2(_0251_ ), .ZN(_0276_ ) );
BUF_X2 _0963_ ( .A(_0276_ ), .Z(_0277_ ) );
INV_X1 _0964_ ( .A(_0277_ ), .ZN(_0278_ ) );
INV_X1 _0965_ ( .A(_0250_ ), .ZN(_0279_ ) );
OAI22_X1 _0966_ ( .A1(_0274_ ), .A2(_0278_ ), .B1(_0279_ ), .B2(_0260_ ), .ZN(_0280_ ) );
AND2_X2 _0967_ ( .A1(_0245_ ), .A2(_0048_ ), .ZN(_0281_ ) );
AND2_X2 _0968_ ( .A1(_0281_ ), .A2(_0249_ ), .ZN(_0282_ ) );
AND2_X1 _0969_ ( .A1(_0282_ ), .A2(_0259_ ), .ZN(_0283_ ) );
BUF_X2 _0970_ ( .A(_0257_ ), .Z(_0284_ ) );
AND2_X1 _0971_ ( .A1(_0284_ ), .A2(_0276_ ), .ZN(_0285_ ) );
AND2_X4 _0972_ ( .A1(_0263_ ), .A2(_0249_ ), .ZN(_0286_ ) );
BUF_X2 _0973_ ( .A(_0286_ ), .Z(_0287_ ) );
BUF_X2 _0974_ ( .A(_0287_ ), .Z(_0288_ ) );
AND2_X1 _0975_ ( .A1(_0288_ ), .A2(_0259_ ), .ZN(_0289_ ) );
NOR4_X1 _0976_ ( .A1(_0280_ ), .A2(_0283_ ), .A3(_0285_ ), .A4(_0289_ ), .ZN(_0290_ ) );
NOR2_X1 _0977_ ( .A1(\inst_o[4] ), .A2(\inst_o[5] ), .ZN(_0291_ ) );
AND2_X2 _0978_ ( .A1(_0251_ ), .A2(_0291_ ), .ZN(_0292_ ) );
AND2_X1 _0979_ ( .A1(_0287_ ), .A2(_0292_ ), .ZN(_0293_ ) );
AND2_X1 _0980_ ( .A1(_0281_ ), .A2(_0269_ ), .ZN(_0294_ ) );
BUF_X2 _0981_ ( .A(_0294_ ), .Z(_0295_ ) );
AND2_X1 _0982_ ( .A1(_0295_ ), .A2(_0292_ ), .ZN(_0296_ ) );
AOI211_X1 _0983_ ( .A(_0293_ ), .B(_0296_ ), .C1(_0282_ ), .C2(_0292_ ), .ZN(_0297_ ) );
NAND2_X1 _0984_ ( .A1(_0282_ ), .A2(_0277_ ), .ZN(_0298_ ) );
NAND2_X1 _0985_ ( .A1(_0295_ ), .A2(_0277_ ), .ZN(_0299_ ) );
NAND2_X1 _0986_ ( .A1(_0288_ ), .A2(_0277_ ), .ZN(_0300_ ) );
AND2_X1 _0987_ ( .A1(_0248_ ), .A2(_0269_ ), .ZN(_0301_ ) );
BUF_X2 _0988_ ( .A(_0301_ ), .Z(_0302_ ) );
NAND2_X1 _0989_ ( .A1(_0302_ ), .A2(_0277_ ), .ZN(_0303_ ) );
AND4_X1 _0990_ ( .A1(_0298_ ), .A2(_0299_ ), .A3(_0300_ ), .A4(_0303_ ), .ZN(_0304_ ) );
AND4_X1 _0991_ ( .A1(_0272_ ), .A2(_0290_ ), .A3(_0297_ ), .A4(_0304_ ), .ZN(_0305_ ) );
AND2_X2 _0992_ ( .A1(_0265_ ), .A2(_0252_ ), .ZN(_0306_ ) );
INV_X1 _0993_ ( .A(_0306_ ), .ZN(_0307_ ) );
INV_X1 _0994_ ( .A(_0301_ ), .ZN(_0308_ ) );
OAI21_X1 _0995_ ( .A(_0249_ ), .B1(_0281_ ), .B2(_0248_ ), .ZN(_0309_ ) );
AOI21_X1 _0996_ ( .A(_0307_ ), .B1(_0308_ ), .B2(_0309_ ), .ZN(_0310_ ) );
AND2_X2 _0997_ ( .A1(_0045_ ), .A2(_0265_ ), .ZN(_0311_ ) );
AND2_X1 _0998_ ( .A1(_0273_ ), .A2(_0311_ ), .ZN(_0312_ ) );
OR2_X1 _0999_ ( .A1(_0310_ ), .A2(_0312_ ), .ZN(_0313_ ) );
NOR2_X1 _1000_ ( .A1(_0295_ ), .A2(_0301_ ), .ZN(_0314_ ) );
AND2_X1 _1001_ ( .A1(_0314_ ), .A2(_0309_ ), .ZN(_0315_ ) );
INV_X1 _1002_ ( .A(\inst_o[6] ), .ZN(_0316_ ) );
NAND3_X1 _1003_ ( .A1(_0316_ ), .A2(_0044_ ), .A3(\inst_o[4] ), .ZN(_0317_ ) );
NOR2_X1 _1004_ ( .A1(_0317_ ), .A2(_0264_ ), .ZN(_0318_ ) );
INV_X1 _1005_ ( .A(_0318_ ), .ZN(_0319_ ) );
NOR2_X1 _1006_ ( .A1(_0315_ ), .A2(_0319_ ), .ZN(_0320_ ) );
AND2_X2 _1007_ ( .A1(_0265_ ), .A2(_0291_ ), .ZN(_0321_ ) );
NOR2_X1 _1008_ ( .A1(_0295_ ), .A2(_0282_ ), .ZN(_0322_ ) );
INV_X1 _1009_ ( .A(_0322_ ), .ZN(_0323_ ) );
AOI211_X1 _1010_ ( .A(_0313_ ), .B(_0320_ ), .C1(_0321_ ), .C2(_0323_ ), .ZN(_0324_ ) );
BUF_X2 _1011_ ( .A(_0253_ ), .Z(_0325_ ) );
OAI21_X1 _1012_ ( .A(_0325_ ), .B1(_0295_ ), .B2(_0288_ ), .ZN(_0326_ ) );
OAI21_X1 _1013_ ( .A(_0325_ ), .B1(_0282_ ), .B2(_0302_ ), .ZN(_0327_ ) );
NAND2_X1 _1014_ ( .A1(_0326_ ), .A2(_0327_ ), .ZN(_0328_ ) );
AND2_X1 _1015_ ( .A1(_0270_ ), .A2(_0259_ ), .ZN(_0329_ ) );
INV_X1 _1016_ ( .A(_0329_ ), .ZN(_0330_ ) );
NAND2_X1 _1017_ ( .A1(_0302_ ), .A2(_0259_ ), .ZN(_0331_ ) );
NAND2_X1 _1018_ ( .A1(_0330_ ), .A2(_0331_ ), .ZN(_0332_ ) );
BUF_X2 _1019_ ( .A(_0270_ ), .Z(_0333_ ) );
AOI211_X1 _1020_ ( .A(_0328_ ), .B(_0332_ ), .C1(_0333_ ), .C2(_0277_ ), .ZN(_0334_ ) );
INV_X1 _1021_ ( .A(_0292_ ), .ZN(_0335_ ) );
AOI21_X1 _1022_ ( .A(_0335_ ), .B1(_0274_ ), .B2(_0258_ ), .ZN(_0336_ ) );
AND2_X1 _1023_ ( .A1(_0333_ ), .A2(_0292_ ), .ZN(_0337_ ) );
NOR2_X1 _1024_ ( .A1(_0336_ ), .A2(_0337_ ), .ZN(_0338_ ) );
AND2_X1 _1025_ ( .A1(_0273_ ), .A2(_0306_ ), .ZN(_0339_ ) );
AND2_X1 _1026_ ( .A1(_0257_ ), .A2(_0306_ ), .ZN(_0340_ ) );
AND2_X1 _1027_ ( .A1(_0270_ ), .A2(_0306_ ), .ZN(_0341_ ) );
AND3_X1 _1028_ ( .A1(_0248_ ), .A2(_0249_ ), .A3(_0292_ ), .ZN(_0342_ ) );
NOR4_X1 _1029_ ( .A1(_0339_ ), .A2(_0340_ ), .A3(_0341_ ), .A4(_0342_ ), .ZN(_0343_ ) );
NAND2_X1 _1030_ ( .A1(_0302_ ), .A2(_0292_ ), .ZN(_0344_ ) );
NAND2_X1 _1031_ ( .A1(_0250_ ), .A2(_0277_ ), .ZN(_0345_ ) );
AND4_X1 _1032_ ( .A1(_0338_ ), .A2(_0343_ ), .A3(_0344_ ), .A4(_0345_ ), .ZN(_0346_ ) );
AND4_X1 _1033_ ( .A1(_0305_ ), .A2(_0324_ ), .A3(_0334_ ), .A4(_0346_ ), .ZN(_0347_ ) );
INV_X1 _1034_ ( .A(_0309_ ), .ZN(_0348_ ) );
OAI21_X1 _1035_ ( .A(_0311_ ), .B1(_0348_ ), .B2(_0302_ ), .ZN(_0349_ ) );
NOR2_X1 _1036_ ( .A1(_0267_ ), .A2(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_ORNOT__Y_A_$_ORNOT__Y_B_$_XOR__A_Y_$_OR__A_1_B ), .ZN(_0350_ ) );
CLKBUF_X2 _1037_ ( .A(_0350_ ), .Z(_0351_ ) );
AND2_X1 _1038_ ( .A1(_0248_ ), .A2(_0351_ ), .ZN(_0352_ ) );
NAND2_X1 _1039_ ( .A1(_0352_ ), .A2(_0311_ ), .ZN(_0353_ ) );
AND2_X1 _1040_ ( .A1(_0349_ ), .A2(_0353_ ), .ZN(_0354_ ) );
BUF_X2 _1041_ ( .A(_0273_ ), .Z(_0355_ ) );
AND2_X1 _1042_ ( .A1(_0355_ ), .A2(_0318_ ), .ZN(_0356_ ) );
AND2_X1 _1043_ ( .A1(_0257_ ), .A2(_0318_ ), .ZN(_0357_ ) );
OR2_X1 _1044_ ( .A1(_0356_ ), .A2(_0357_ ), .ZN(_0358_ ) );
OR2_X1 _1045_ ( .A1(_0295_ ), .A2(_0288_ ), .ZN(_0359_ ) );
AND2_X1 _1046_ ( .A1(_0359_ ), .A2(_0306_ ), .ZN(_0360_ ) );
INV_X1 _1047_ ( .A(_0311_ ), .ZN(_0361_ ) );
INV_X1 _1048_ ( .A(_0333_ ), .ZN(_0362_ ) );
AOI21_X1 _1049_ ( .A(_0361_ ), .B1(_0258_ ), .B2(_0362_ ), .ZN(_0363_ ) );
INV_X1 _1050_ ( .A(_0295_ ), .ZN(_0364_ ) );
INV_X1 _1051_ ( .A(_0288_ ), .ZN(_0365_ ) );
AOI21_X1 _1052_ ( .A(_0361_ ), .B1(_0364_ ), .B2(_0365_ ), .ZN(_0366_ ) );
NOR4_X1 _1053_ ( .A1(_0358_ ), .A2(_0360_ ), .A3(_0363_ ), .A4(_0366_ ), .ZN(_0367_ ) );
OAI21_X1 _1054_ ( .A(_0318_ ), .B1(_0333_ ), .B2(_0288_ ), .ZN(_0368_ ) );
BUF_X2 _1055_ ( .A(_0255_ ), .Z(_0369_ ) );
BUF_X4 _1056_ ( .A(_0249_ ), .Z(_0370_ ) );
BUF_X4 _1057_ ( .A(_0269_ ), .Z(_0371_ ) );
OAI211_X1 _1058_ ( .A(_0369_ ), .B(_0321_ ), .C1(_0370_ ), .C2(_0371_ ), .ZN(_0372_ ) );
AND2_X1 _1059_ ( .A1(_0368_ ), .A2(_0372_ ), .ZN(_0373_ ) );
BUF_X4 _1060_ ( .A(_0263_ ), .Z(_0374_ ) );
BUF_X4 _1061_ ( .A(_0374_ ), .Z(_0375_ ) );
OAI221_X1 _1062_ ( .A(_0321_ ), .B1(_0370_ ), .B2(_0371_ ), .C1(_0248_ ), .C2(_0375_ ), .ZN(_0376_ ) );
AND4_X1 _1063_ ( .A1(_0354_ ), .A2(_0367_ ), .A3(_0373_ ), .A4(_0376_ ), .ZN(_0377_ ) );
AOI21_X1 _1064_ ( .A(reset ), .B1(_0347_ ), .B2(_0377_ ), .ZN(_0036_ ) );
NOR2_X1 _1065_ ( .A1(_0333_ ), .A2(_0288_ ), .ZN(_0378_ ) );
AOI21_X1 _1066_ ( .A(_0278_ ), .B1(_0315_ ), .B2(_0378_ ), .ZN(_0379_ ) );
AND2_X1 _1067_ ( .A1(_0355_ ), .A2(_0277_ ), .ZN(_0380_ ) );
OR2_X1 _1068_ ( .A1(_0380_ ), .A2(_0285_ ), .ZN(_0381_ ) );
NOR2_X1 _1069_ ( .A1(_0379_ ), .A2(_0381_ ), .ZN(_0382_ ) );
NOR2_X1 _1070_ ( .A1(_0316_ ), .A2(\inst_o[7] ), .ZN(_0383_ ) );
AND2_X1 _1071_ ( .A1(_0383_ ), .A2(_0252_ ), .ZN(_0384_ ) );
BUF_X2 _1072_ ( .A(_0384_ ), .Z(_0385_ ) );
AND2_X1 _1073_ ( .A1(_0273_ ), .A2(_0385_ ), .ZN(_0386_ ) );
AND2_X1 _1074_ ( .A1(_0288_ ), .A2(_0325_ ), .ZN(_0387_ ) );
NOR4_X1 _1075_ ( .A1(_0262_ ), .A2(_0386_ ), .A3(_0387_ ), .A4(_0271_ ), .ZN(_0388_ ) );
INV_X1 _1076_ ( .A(_0325_ ), .ZN(_0389_ ) );
NOR2_X1 _1077_ ( .A1(_0322_ ), .A2(_0389_ ), .ZN(_0390_ ) );
INV_X1 _1078_ ( .A(_0390_ ), .ZN(_0391_ ) );
NAND2_X1 _1079_ ( .A1(_0388_ ), .A2(_0391_ ), .ZN(_0392_ ) );
AOI21_X1 _1080_ ( .A(_0335_ ), .B1(_0315_ ), .B2(_0365_ ), .ZN(_0393_ ) );
NOR2_X1 _1081_ ( .A1(_0392_ ), .A2(_0393_ ), .ZN(_0394_ ) );
INV_X1 _1082_ ( .A(_0378_ ), .ZN(_0395_ ) );
AND2_X1 _1083_ ( .A1(_0045_ ), .A2(_0383_ ), .ZN(_0396_ ) );
BUF_X2 _1084_ ( .A(_0396_ ), .Z(_0397_ ) );
AND2_X1 _1085_ ( .A1(_0383_ ), .A2(_0291_ ), .ZN(_0398_ ) );
BUF_X2 _1086_ ( .A(_0398_ ), .Z(_0399_ ) );
OAI21_X1 _1087_ ( .A(_0395_ ), .B1(_0397_ ), .B2(_0399_ ), .ZN(_0400_ ) );
AND2_X1 _1088_ ( .A1(_0275_ ), .A2(_0383_ ), .ZN(_0401_ ) );
INV_X1 _1089_ ( .A(_0401_ ), .ZN(_0402_ ) );
AOI21_X1 _1090_ ( .A(_0402_ ), .B1(_0308_ ), .B2(_0279_ ), .ZN(_0403_ ) );
BUF_X2 _1091_ ( .A(_0401_ ), .Z(_0404_ ) );
AOI21_X1 _1092_ ( .A(_0403_ ), .B1(_0323_ ), .B2(_0404_ ), .ZN(_0405_ ) );
AND4_X1 _1093_ ( .A1(_0382_ ), .A2(_0394_ ), .A3(_0400_ ), .A4(_0405_ ), .ZN(_0406_ ) );
AND2_X1 _1094_ ( .A1(_0257_ ), .A2(_0396_ ), .ZN(_0407_ ) );
AND2_X1 _1095_ ( .A1(_0282_ ), .A2(_0397_ ), .ZN(_0408_ ) );
NOR2_X1 _1096_ ( .A1(_0407_ ), .A2(_0408_ ), .ZN(_0409_ ) );
AND2_X1 _1097_ ( .A1(_0322_ ), .A2(_0258_ ), .ZN(_0410_ ) );
AND2_X1 _1098_ ( .A1(_0410_ ), .A2(_0274_ ), .ZN(_0411_ ) );
INV_X1 _1099_ ( .A(_0398_ ), .ZN(_0412_ ) );
OAI21_X1 _1100_ ( .A(_0409_ ), .B1(_0411_ ), .B2(_0412_ ), .ZN(_0413_ ) );
NOR3_X1 _1101_ ( .A1(_0284_ ), .A2(_0333_ ), .A3(_0288_ ), .ZN(_0414_ ) );
INV_X1 _1102_ ( .A(_0384_ ), .ZN(_0415_ ) );
OR2_X1 _1103_ ( .A1(_0414_ ), .A2(_0415_ ), .ZN(_0416_ ) );
OAI21_X1 _1104_ ( .A(_0404_ ), .B1(_0355_ ), .B2(_0284_ ), .ZN(_0417_ ) );
OAI211_X1 _1105_ ( .A(_0375_ ), .B(_0404_ ), .C1(_0370_ ), .C2(_0269_ ), .ZN(_0418_ ) );
AND2_X1 _1106_ ( .A1(_0417_ ), .A2(_0418_ ), .ZN(_0419_ ) );
OAI211_X1 _1107_ ( .A(_0416_ ), .B(_0419_ ), .C1(_0315_ ), .C2(_0415_ ), .ZN(_0420_ ) );
NAND2_X1 _1108_ ( .A1(_0302_ ), .A2(_0396_ ), .ZN(_0421_ ) );
NAND2_X1 _1109_ ( .A1(_0250_ ), .A2(_0397_ ), .ZN(_0422_ ) );
OAI21_X1 _1110_ ( .A(_0259_ ), .B1(_0284_ ), .B2(_0333_ ), .ZN(_0423_ ) );
NAND4_X1 _1111_ ( .A1(_0338_ ), .A2(_0421_ ), .A3(_0422_ ), .A4(_0423_ ), .ZN(_0424_ ) );
NOR2_X1 _1112_ ( .A1(_0283_ ), .A2(_0289_ ), .ZN(_0425_ ) );
OAI221_X1 _1113_ ( .A(_0248_ ), .B1(_0371_ ), .B2(_0370_ ), .C1(_0325_ ), .C2(_0399_ ), .ZN(_0426_ ) );
NOR2_X1 _1114_ ( .A1(_0302_ ), .A2(_0250_ ), .ZN(_0427_ ) );
OAI211_X1 _1115_ ( .A(_0425_ ), .B(_0426_ ), .C1(_0260_ ), .C2(_0427_ ), .ZN(_0428_ ) );
NOR4_X1 _1116_ ( .A1(_0413_ ), .A2(_0420_ ), .A3(_0424_ ), .A4(_0428_ ), .ZN(_0429_ ) );
AOI21_X1 _1117_ ( .A(reset ), .B1(_0406_ ), .B2(_0429_ ), .ZN(_0037_ ) );
OR2_X1 _1118_ ( .A1(_0283_ ), .A2(_0339_ ), .ZN(_0430_ ) );
OR4_X1 _1119_ ( .A1(_0289_ ), .A2(_0430_ ), .A3(_0261_ ), .A4(_0329_ ), .ZN(_0431_ ) );
AND2_X1 _1120_ ( .A1(_0250_ ), .A2(_0397_ ), .ZN(_0432_ ) );
NOR2_X1 _1121_ ( .A1(_0262_ ), .A2(_0386_ ), .ZN(_0433_ ) );
OAI221_X1 _1122_ ( .A(_0433_ ), .B1(_0362_ ), .B2(_0389_ ), .C1(_0260_ ), .C2(_0427_ ), .ZN(_0434_ ) );
NOR4_X1 _1123_ ( .A1(_0431_ ), .A2(_0328_ ), .A3(_0432_ ), .A4(_0434_ ), .ZN(_0435_ ) );
NOR2_X1 _1124_ ( .A1(\inst_o[6] ), .A2(\inst_o[7] ), .ZN(_0436_ ) );
AND2_X1 _1125_ ( .A1(_0252_ ), .A2(_0436_ ), .ZN(_0437_ ) );
BUF_X2 _1126_ ( .A(_0437_ ), .Z(_0438_ ) );
OAI21_X1 _1127_ ( .A(_0438_ ), .B1(_0284_ ), .B2(_0333_ ), .ZN(_0439_ ) );
NAND2_X1 _1128_ ( .A1(_0295_ ), .A2(_0438_ ), .ZN(_0440_ ) );
INV_X1 _1129_ ( .A(_0438_ ), .ZN(_0441_ ) );
OAI211_X1 _1130_ ( .A(_0439_ ), .B(_0440_ ), .C1(_0365_ ), .C2(_0441_ ), .ZN(_0442_ ) );
AND2_X1 _1131_ ( .A1(_0045_ ), .A2(_0436_ ), .ZN(_0443_ ) );
BUF_X2 _1132_ ( .A(_0443_ ), .Z(_0444_ ) );
NAND2_X1 _1133_ ( .A1(_0333_ ), .A2(_0444_ ), .ZN(_0445_ ) );
NAND2_X1 _1134_ ( .A1(_0286_ ), .A2(_0444_ ), .ZN(_0446_ ) );
INV_X1 _1135_ ( .A(_0444_ ), .ZN(_0447_ ) );
OAI211_X1 _1136_ ( .A(_0445_ ), .B(_0446_ ), .C1(_0364_ ), .C2(_0447_ ), .ZN(_0448_ ) );
AOI21_X1 _1137_ ( .A(_0447_ ), .B1(_0308_ ), .B2(_0309_ ), .ZN(_0449_ ) );
AOI21_X1 _1138_ ( .A(_0415_ ), .B1(_0308_ ), .B2(_0309_ ), .ZN(_0450_ ) );
NOR4_X1 _1139_ ( .A1(_0442_ ), .A2(_0448_ ), .A3(_0449_ ), .A4(_0450_ ), .ZN(_0451_ ) );
OAI22_X1 _1140_ ( .A1(_0274_ ), .A2(_0447_ ), .B1(_0279_ ), .B2(_0441_ ), .ZN(_0452_ ) );
AND2_X1 _1141_ ( .A1(_0256_ ), .A2(_0444_ ), .ZN(_0453_ ) );
AND2_X1 _1142_ ( .A1(_0282_ ), .A2(_0438_ ), .ZN(_0454_ ) );
AND2_X1 _1143_ ( .A1(_0302_ ), .A2(_0438_ ), .ZN(_0455_ ) );
NOR4_X1 _1144_ ( .A1(_0452_ ), .A2(_0453_ ), .A3(_0454_ ), .A4(_0455_ ), .ZN(_0456_ ) );
AOI21_X1 _1145_ ( .A(_0408_ ), .B1(_0395_ ), .B2(_0397_ ), .ZN(_0457_ ) );
OAI21_X1 _1146_ ( .A(_0397_ ), .B1(_0284_ ), .B2(_0302_ ), .ZN(_0458_ ) );
AOI22_X1 _1147_ ( .A1(_0355_ ), .A2(_0438_ ), .B1(_0295_ ), .B2(_0385_ ), .ZN(_0459_ ) );
AND4_X1 _1148_ ( .A1(_0416_ ), .A2(_0457_ ), .A3(_0458_ ), .A4(_0459_ ), .ZN(_0460_ ) );
AND4_X1 _1149_ ( .A1(_0435_ ), .A2(_0451_ ), .A3(_0456_ ), .A4(_0460_ ), .ZN(_0461_ ) );
OR3_X1 _1150_ ( .A1(_0360_ ), .A2(_0341_ ), .A3(_0340_ ), .ZN(_0462_ ) );
NAND2_X1 _1151_ ( .A1(_0287_ ), .A2(_0311_ ), .ZN(_0463_ ) );
OAI211_X1 _1152_ ( .A(_0354_ ), .B(_0463_ ), .C1(_0361_ ), .C2(_0364_ ), .ZN(_0464_ ) );
NOR4_X1 _1153_ ( .A1(_0462_ ), .A2(_0464_ ), .A3(_0313_ ), .A4(_0363_ ), .ZN(_0465_ ) );
AOI21_X1 _1154_ ( .A(reset ), .B1(_0461_ ), .B2(_0465_ ), .ZN(_0038_ ) );
NOR2_X1 _1155_ ( .A1(_0317_ ), .A2(\inst_o[7] ), .ZN(_0466_ ) );
BUF_X2 _1156_ ( .A(_0466_ ), .Z(_0467_ ) );
AND2_X1 _1157_ ( .A1(_0256_ ), .A2(_0467_ ), .ZN(_0468_ ) );
NOR3_X1 _1158_ ( .A1(_0339_ ), .A2(_0340_ ), .A3(_0468_ ), .ZN(_0469_ ) );
NOR2_X1 _1159_ ( .A1(_0356_ ), .A2(_0357_ ), .ZN(_0470_ ) );
INV_X1 _1160_ ( .A(_0314_ ), .ZN(_0471_ ) );
OAI22_X1 _1161_ ( .A1(_0471_ ), .A2(_0348_ ), .B1(_0318_ ), .B2(_0385_ ), .ZN(_0472_ ) );
AND4_X1 _1162_ ( .A1(_0368_ ), .A2(_0469_ ), .A3(_0470_ ), .A4(_0472_ ), .ZN(_0473_ ) );
OAI22_X1 _1163_ ( .A1(_0471_ ), .A2(_0348_ ), .B1(_0306_ ), .B2(_0438_ ), .ZN(_0474_ ) );
OAI21_X1 _1164_ ( .A(_0467_ ), .B1(_0471_ ), .B2(_0348_ ), .ZN(_0475_ ) );
AND3_X1 _1165_ ( .A1(_0474_ ), .A2(_0475_ ), .A3(_0419_ ), .ZN(_0476_ ) );
OAI21_X1 _1166_ ( .A(_0395_ ), .B1(_0306_ ), .B2(_0467_ ), .ZN(_0477_ ) );
OR2_X1 _1167_ ( .A1(_0322_ ), .A2(_0402_ ), .ZN(_0478_ ) );
OAI221_X1 _1168_ ( .A(_0248_ ), .B1(_0371_ ), .B2(_0370_ ), .C1(_0325_ ), .C2(_0404_ ), .ZN(_0479_ ) );
AND3_X1 _1169_ ( .A1(_0477_ ), .A2(_0478_ ), .A3(_0479_ ), .ZN(_0480_ ) );
AND4_X1 _1170_ ( .A1(_0382_ ), .A2(_0473_ ), .A3(_0476_ ), .A4(_0480_ ), .ZN(_0481_ ) );
NAND2_X1 _1171_ ( .A1(_0355_ ), .A2(_0438_ ), .ZN(_0482_ ) );
NAND2_X1 _1172_ ( .A1(_0416_ ), .A2(_0482_ ), .ZN(_0483_ ) );
AND2_X1 _1173_ ( .A1(_0355_ ), .A2(_0467_ ), .ZN(_0484_ ) );
AND2_X1 _1174_ ( .A1(_0286_ ), .A2(_0437_ ), .ZN(_0485_ ) );
NOR2_X1 _1175_ ( .A1(_0484_ ), .A2(_0485_ ), .ZN(_0486_ ) );
NAND2_X1 _1176_ ( .A1(_0486_ ), .A2(_0439_ ), .ZN(_0487_ ) );
NOR3_X1 _1177_ ( .A1(_0392_ ), .A2(_0483_ ), .A3(_0487_ ), .ZN(_0488_ ) );
AOI21_X1 _1178_ ( .A(reset ), .B1(_0481_ ), .B2(_0488_ ), .ZN(_0039_ ) );
NOR2_X1 _1179_ ( .A1(_0358_ ), .A2(_0381_ ), .ZN(_0489_ ) );
OAI211_X1 _1180_ ( .A(_0489_ ), .B(_0373_ ), .C1(_0361_ ), .C2(_0414_ ), .ZN(_0490_ ) );
NOR4_X1 _1181_ ( .A1(_0312_ ), .A2(_0339_ ), .A3(_0340_ ), .A4(_0337_ ), .ZN(_0491_ ) );
AND2_X1 _1182_ ( .A1(_0273_ ), .A2(_0399_ ), .ZN(_0492_ ) );
AND2_X1 _1183_ ( .A1(_0256_ ), .A2(_0398_ ), .ZN(_0493_ ) );
AND2_X1 _1184_ ( .A1(_0291_ ), .A2(_0436_ ), .ZN(_0494_ ) );
BUF_X2 _1185_ ( .A(_0494_ ), .Z(_0495_ ) );
AND2_X1 _1186_ ( .A1(_0355_ ), .A2(_0495_ ), .ZN(_0496_ ) );
NOR4_X1 _1187_ ( .A1(_0492_ ), .A2(_0493_ ), .A3(_0496_ ), .A4(_0293_ ), .ZN(_0497_ ) );
AND2_X2 _1188_ ( .A1(_0286_ ), .A2(_0495_ ), .ZN(_0498_ ) );
NOR4_X1 _1189_ ( .A1(_0386_ ), .A2(_0407_ ), .A3(_0468_ ), .A4(_0498_ ), .ZN(_0499_ ) );
NOR3_X1 _1190_ ( .A1(_0336_ ), .A2(_0262_ ), .A3(_0271_ ), .ZN(_0500_ ) );
NAND4_X1 _1191_ ( .A1(_0491_ ), .A2(_0497_ ), .A3(_0499_ ), .A4(_0500_ ), .ZN(_0501_ ) );
AOI21_X1 _1192_ ( .A(_0378_ ), .B1(_0260_ ), .B2(_0447_ ), .ZN(_0502_ ) );
AND2_X1 _1193_ ( .A1(_0273_ ), .A2(_0444_ ), .ZN(_0503_ ) );
NOR3_X1 _1194_ ( .A1(_0502_ ), .A2(_0503_ ), .A3(_0453_ ), .ZN(_0504_ ) );
OAI221_X1 _1195_ ( .A(_0375_ ), .B1(_0371_ ), .B2(_0370_ ), .C1(_0321_ ), .C2(_0277_ ), .ZN(_0505_ ) );
NAND4_X1 _1196_ ( .A1(_0504_ ), .A2(_0400_ ), .A3(_0419_ ), .A4(_0505_ ), .ZN(_0506_ ) );
NOR3_X1 _1197_ ( .A1(_0490_ ), .A2(_0501_ ), .A3(_0506_ ), .ZN(_0507_ ) );
NAND2_X1 _1198_ ( .A1(_0256_ ), .A2(_0495_ ), .ZN(_0508_ ) );
NAND2_X1 _1199_ ( .A1(_0270_ ), .A2(_0495_ ), .ZN(_0509_ ) );
NAND3_X1 _1200_ ( .A1(_0477_ ), .A2(_0508_ ), .A3(_0509_ ), .ZN(_0510_ ) );
NAND2_X1 _1201_ ( .A1(_0288_ ), .A2(_0325_ ), .ZN(_0511_ ) );
OAI21_X1 _1202_ ( .A(_0511_ ), .B1(_0258_ ), .B2(_0260_ ), .ZN(_0512_ ) );
NOR4_X1 _1203_ ( .A1(_0483_ ), .A2(_0510_ ), .A3(_0487_ ), .A4(_0512_ ), .ZN(_0513_ ) );
AOI21_X1 _1204_ ( .A(reset ), .B1(_0507_ ), .B2(_0513_ ), .ZN(_0040_ ) );
INV_X1 _1205_ ( .A(_0262_ ), .ZN(_0514_ ) );
OAI21_X1 _1206_ ( .A(_0399_ ), .B1(_0282_ ), .B2(_0295_ ), .ZN(_0515_ ) );
AND2_X1 _1207_ ( .A1(_0251_ ), .A2(_0044_ ), .ZN(_0516_ ) );
OAI221_X1 _1208_ ( .A(_0516_ ), .B1(_0370_ ), .B2(_0371_ ), .C1(_0281_ ), .C2(_0369_ ), .ZN(_0517_ ) );
AND3_X1 _1209_ ( .A1(_0514_ ), .A2(_0515_ ), .A3(_0517_ ), .ZN(_0518_ ) );
OAI21_X1 _1210_ ( .A(_0385_ ), .B1(_0323_ ), .B2(_0284_ ), .ZN(_0519_ ) );
OAI221_X1 _1211_ ( .A(_0444_ ), .B1(_0370_ ), .B2(_0371_ ), .C1(_0281_ ), .C2(_0369_ ), .ZN(_0520_ ) );
AND2_X1 _1212_ ( .A1(_0519_ ), .A2(_0520_ ), .ZN(_0521_ ) );
AND2_X1 _1213_ ( .A1(_0284_ ), .A2(_0259_ ), .ZN(_0522_ ) );
NOR4_X1 _1214_ ( .A1(_0390_ ), .A2(_0283_ ), .A3(_0522_ ), .A4(_0386_ ), .ZN(_0523_ ) );
OAI221_X1 _1215_ ( .A(_0265_ ), .B1(_0370_ ), .B2(_0371_ ), .C1(_0281_ ), .C2(_0369_ ), .ZN(_0524_ ) );
AND4_X1 _1216_ ( .A1(_0518_ ), .A2(_0521_ ), .A3(_0523_ ), .A4(_0524_ ), .ZN(_0525_ ) );
OAI22_X1 _1217_ ( .A1(_0323_ ), .A2(_0284_ ), .B1(_0438_ ), .B2(_0467_ ), .ZN(_0526_ ) );
OAI221_X1 _1218_ ( .A(_0369_ ), .B1(_0370_ ), .B2(_0269_ ), .C1(_0399_ ), .C2(_0404_ ), .ZN(_0527_ ) );
AND4_X1 _1219_ ( .A1(_0478_ ), .A2(_0409_ ), .A3(_0482_ ), .A4(_0527_ ), .ZN(_0528_ ) );
OAI21_X1 _1220_ ( .A(_0495_ ), .B1(_0323_ ), .B2(_0284_ ), .ZN(_0529_ ) );
OAI211_X1 _1221_ ( .A(_0369_ ), .B(_0371_ ), .C1(_0467_ ), .C2(_0495_ ), .ZN(_0530_ ) );
AND4_X1 _1222_ ( .A1(_0526_ ), .A2(_0528_ ), .A3(_0529_ ), .A4(_0530_ ), .ZN(_0531_ ) );
AOI21_X1 _1223_ ( .A(reset ), .B1(_0525_ ), .B2(_0531_ ), .ZN(_0041_ ) );
INV_X1 _1224_ ( .A(_0289_ ), .ZN(_0532_ ) );
AND2_X1 _1225_ ( .A1(_0257_ ), .A2(_0292_ ), .ZN(_0533_ ) );
INV_X1 _1226_ ( .A(_0293_ ), .ZN(_0534_ ) );
AND2_X1 _1227_ ( .A1(_0287_ ), .A2(_0306_ ), .ZN(_0535_ ) );
INV_X1 _1228_ ( .A(_0535_ ), .ZN(_0536_ ) );
AND2_X1 _1229_ ( .A1(_0257_ ), .A2(_0311_ ), .ZN(_0537_ ) );
NAND2_X1 _1230_ ( .A1(_0287_ ), .A2(_0318_ ), .ZN(_0538_ ) );
AND2_X1 _1231_ ( .A1(_0257_ ), .A2(_0321_ ), .ZN(_0539_ ) );
NAND2_X1 _1232_ ( .A1(_0287_ ), .A2(_0321_ ), .ZN(_0540_ ) );
AND2_X1 _1233_ ( .A1(_0257_ ), .A2(_0385_ ), .ZN(_0541_ ) );
NAND2_X1 _1234_ ( .A1(_0287_ ), .A2(_0385_ ), .ZN(_0542_ ) );
NAND2_X1 _1235_ ( .A1(_0287_ ), .A2(_0396_ ), .ZN(_0543_ ) );
AND2_X1 _1236_ ( .A1(_0256_ ), .A2(_0401_ ), .ZN(_0544_ ) );
NAND2_X1 _1237_ ( .A1(_0287_ ), .A2(_0404_ ), .ZN(_0545_ ) );
NAND2_X1 _1238_ ( .A1(_0287_ ), .A2(_0399_ ), .ZN(_0546_ ) );
AND2_X1 _1239_ ( .A1(_0256_ ), .A2(_0437_ ), .ZN(_0547_ ) );
INV_X1 _1240_ ( .A(_0485_ ), .ZN(_0548_ ) );
NAND3_X1 _1241_ ( .A1(_0255_ ), .A2(_0351_ ), .A3(_0467_ ), .ZN(_0549_ ) );
AND3_X1 _1242_ ( .A1(_0281_ ), .A2(_0351_ ), .A3(_0443_ ), .ZN(_0550_ ) );
AOI221_X4 _1243_ ( .A(_0550_ ), .B1(_0352_ ), .B2(_0444_ ), .C1(_0273_ ), .C2(_0467_ ), .ZN(_0551_ ) );
AND3_X1 _1244_ ( .A1(_0374_ ), .A2(_0351_ ), .A3(_0466_ ), .ZN(_0552_ ) );
NAND3_X1 _1245_ ( .A1(_0374_ ), .A2(_0350_ ), .A3(_0495_ ), .ZN(_0553_ ) );
OAI221_X1 _1246_ ( .A(_0495_ ), .B1(_0350_ ), .B2(_0269_ ), .C1(_0281_ ), .C2(_0248_ ), .ZN(_0554_ ) );
OAI211_X1 _1247_ ( .A(_0509_ ), .B(_0553_ ), .C1(_0498_ ), .C2(_0554_ ), .ZN(_0555_ ) );
NAND2_X1 _1248_ ( .A1(_0555_ ), .A2(_0508_ ), .ZN(_0556_ ) );
OAI21_X1 _1249_ ( .A(_0466_ ), .B1(_0294_ ), .B2(_0301_ ), .ZN(_0557_ ) );
NAND3_X1 _1250_ ( .A1(_0255_ ), .A2(_0351_ ), .A3(_0495_ ), .ZN(_0558_ ) );
AND3_X1 _1251_ ( .A1(_0247_ ), .A2(_0350_ ), .A3(_0466_ ), .ZN(_0559_ ) );
AND2_X1 _1252_ ( .A1(_0281_ ), .A2(_0350_ ), .ZN(_0560_ ) );
AOI221_X2 _1253_ ( .A(_0559_ ), .B1(_0273_ ), .B2(_0494_ ), .C1(_0466_ ), .C2(_0560_ ), .ZN(_0561_ ) );
NAND4_X1 _1254_ ( .A1(_0556_ ), .A2(_0557_ ), .A3(_0558_ ), .A4(_0561_ ), .ZN(_0562_ ) );
NAND2_X1 _1255_ ( .A1(_0286_ ), .A2(_0466_ ), .ZN(_0563_ ) );
AOI221_X1 _1256_ ( .A(_0552_ ), .B1(_0270_ ), .B2(_0467_ ), .C1(_0562_ ), .C2(_0563_ ), .ZN(_0564_ ) );
OAI211_X1 _1257_ ( .A(_0549_ ), .B(_0551_ ), .C1(_0564_ ), .C2(_0468_ ), .ZN(_0565_ ) );
AOI21_X1 _1258_ ( .A(_0447_ ), .B1(_0364_ ), .B2(_0308_ ), .ZN(_0566_ ) );
OAI21_X1 _1259_ ( .A(_0446_ ), .B1(_0565_ ), .B2(_0566_ ), .ZN(_0567_ ) );
NAND3_X1 _1260_ ( .A1(_0374_ ), .A2(_0268_ ), .A3(_0444_ ), .ZN(_0568_ ) );
AOI21_X1 _1261_ ( .A(_0453_ ), .B1(_0567_ ), .B2(_0568_ ), .ZN(_0569_ ) );
AND2_X1 _1262_ ( .A1(_0437_ ), .A2(_0268_ ), .ZN(_0570_ ) );
AND3_X1 _1263_ ( .A1(_0245_ ), .A2(_0048_ ), .A3(_0570_ ), .ZN(_0571_ ) );
INV_X1 _1264_ ( .A(_0570_ ), .ZN(_0572_ ) );
NOR3_X1 _1265_ ( .A1(_0245_ ), .A2(_0246_ ), .A3(_0572_ ), .ZN(_0573_ ) );
AND3_X1 _1266_ ( .A1(_0255_ ), .A2(_0351_ ), .A3(_0444_ ), .ZN(_0574_ ) );
OR4_X1 _1267_ ( .A1(_0571_ ), .A2(_0503_ ), .A3(_0573_ ), .A4(_0574_ ), .ZN(_0575_ ) );
OAI21_X1 _1268_ ( .A(_0548_ ), .B1(_0569_ ), .B2(_0575_ ), .ZN(_0576_ ) );
NOR3_X1 _1269_ ( .A1(_0245_ ), .A2(_0048_ ), .A3(_0572_ ), .ZN(_0577_ ) );
INV_X1 _1270_ ( .A(_0577_ ), .ZN(_0578_ ) );
AOI21_X1 _1271_ ( .A(_0547_ ), .B1(_0576_ ), .B2(_0578_ ), .ZN(_0579_ ) );
INV_X1 _1272_ ( .A(_0243_ ), .ZN(_0580_ ) );
NAND4_X1 _1273_ ( .A1(_0580_ ), .A2(\inst_o[2] ), .A3(_0246_ ), .A4(_0570_ ), .ZN(_0581_ ) );
OR2_X1 _1274_ ( .A1(_0560_ ), .A2(_0352_ ), .ZN(_0582_ ) );
NOR2_X1 _1275_ ( .A1(_0471_ ), .A2(_0582_ ), .ZN(_0583_ ) );
OAI21_X1 _1276_ ( .A(_0581_ ), .B1(_0583_ ), .B2(_0412_ ), .ZN(_0584_ ) );
OAI21_X1 _1277_ ( .A(_0546_ ), .B1(_0579_ ), .B2(_0584_ ), .ZN(_0585_ ) );
NAND3_X1 _1278_ ( .A1(_0374_ ), .A2(_0268_ ), .A3(_0399_ ), .ZN(_0586_ ) );
AOI21_X1 _1279_ ( .A(_0493_ ), .B1(_0585_ ), .B2(_0586_ ), .ZN(_0587_ ) );
NAND3_X1 _1280_ ( .A1(_0255_ ), .A2(_0351_ ), .A3(_0399_ ), .ZN(_0588_ ) );
OAI221_X1 _1281_ ( .A(_0588_ ), .B1(_0274_ ), .B2(_0412_ ), .C1(_0583_ ), .C2(_0402_ ), .ZN(_0589_ ) );
OAI21_X1 _1282_ ( .A(_0545_ ), .B1(_0587_ ), .B2(_0589_ ), .ZN(_0590_ ) );
NAND3_X1 _1283_ ( .A1(_0374_ ), .A2(_0268_ ), .A3(_0404_ ), .ZN(_0591_ ) );
AOI21_X1 _1284_ ( .A(_0544_ ), .B1(_0590_ ), .B2(_0591_ ), .ZN(_0592_ ) );
OAI21_X1 _1285_ ( .A(_0396_ ), .B1(_0560_ ), .B2(_0352_ ), .ZN(_0593_ ) );
NAND2_X1 _1286_ ( .A1(_0369_ ), .A2(_0268_ ), .ZN(_0594_ ) );
OAI211_X1 _1287_ ( .A(_0593_ ), .B(_0421_ ), .C1(_0402_ ), .C2(_0594_ ), .ZN(_0595_ ) );
OAI21_X1 _1288_ ( .A(_0543_ ), .B1(_0592_ ), .B2(_0595_ ), .ZN(_0596_ ) );
NAND3_X1 _1289_ ( .A1(_0374_ ), .A2(_0268_ ), .A3(_0397_ ), .ZN(_0597_ ) );
AOI21_X1 _1290_ ( .A(_0407_ ), .B1(_0596_ ), .B2(_0597_ ), .ZN(_0598_ ) );
NAND3_X1 _1291_ ( .A1(_0369_ ), .A2(_0351_ ), .A3(_0397_ ), .ZN(_0599_ ) );
OAI21_X1 _1292_ ( .A(_0599_ ), .B1(_0583_ ), .B2(_0415_ ), .ZN(_0600_ ) );
OAI21_X1 _1293_ ( .A(_0542_ ), .B1(_0598_ ), .B2(_0600_ ), .ZN(_0601_ ) );
BUF_X4 _1294_ ( .A(_0268_ ), .Z(_0602_ ) );
NAND3_X1 _1295_ ( .A1(_0374_ ), .A2(_0602_ ), .A3(_0385_ ), .ZN(_0603_ ) );
AOI21_X1 _1296_ ( .A(_0541_ ), .B1(_0601_ ), .B2(_0603_ ), .ZN(_0604_ ) );
INV_X1 _1297_ ( .A(_0321_ ), .ZN(_0605_ ) );
OAI22_X1 _1298_ ( .A1(_0583_ ), .A2(_0605_ ), .B1(_0415_ ), .B2(_0594_ ), .ZN(_0606_ ) );
OAI21_X1 _1299_ ( .A(_0540_ ), .B1(_0604_ ), .B2(_0606_ ), .ZN(_0607_ ) );
NAND3_X1 _1300_ ( .A1(_0374_ ), .A2(_0602_ ), .A3(_0321_ ), .ZN(_0608_ ) );
AOI21_X1 _1301_ ( .A(_0539_ ), .B1(_0607_ ), .B2(_0608_ ), .ZN(_0609_ ) );
OAI22_X1 _1302_ ( .A1(_0583_ ), .A2(_0319_ ), .B1(_0605_ ), .B2(_0594_ ), .ZN(_0610_ ) );
OAI21_X1 _1303_ ( .A(_0538_ ), .B1(_0609_ ), .B2(_0610_ ), .ZN(_0611_ ) );
NAND3_X1 _1304_ ( .A1(_0374_ ), .A2(_0602_ ), .A3(_0318_ ), .ZN(_0612_ ) );
AOI21_X1 _1305_ ( .A(_0357_ ), .B1(_0611_ ), .B2(_0612_ ), .ZN(_0613_ ) );
AOI22_X1 _1306_ ( .A1(_0281_ ), .A2(_0602_ ), .B1(_0248_ ), .B2(_0269_ ), .ZN(_0614_ ) );
OAI221_X1 _1307_ ( .A(_0353_ ), .B1(_0319_ ), .B2(_0594_ ), .C1(_0614_ ), .C2(_0361_ ), .ZN(_0615_ ) );
OAI21_X1 _1308_ ( .A(_0463_ ), .B1(_0613_ ), .B2(_0615_ ), .ZN(_0616_ ) );
NAND3_X1 _1309_ ( .A1(_0375_ ), .A2(_0602_ ), .A3(_0311_ ), .ZN(_0617_ ) );
AOI21_X1 _1310_ ( .A(_0537_ ), .B1(_0616_ ), .B2(_0617_ ), .ZN(_0618_ ) );
OAI22_X1 _1311_ ( .A1(_0583_ ), .A2(_0307_ ), .B1(_0361_ ), .B2(_0594_ ), .ZN(_0619_ ) );
OAI21_X1 _1312_ ( .A(_0536_ ), .B1(_0618_ ), .B2(_0619_ ), .ZN(_0620_ ) );
NAND3_X1 _1313_ ( .A1(_0375_ ), .A2(_0602_ ), .A3(_0306_ ), .ZN(_0621_ ) );
AOI21_X1 _1314_ ( .A(_0340_ ), .B1(_0620_ ), .B2(_0621_ ), .ZN(_0622_ ) );
OAI22_X1 _1315_ ( .A1(_0583_ ), .A2(_0335_ ), .B1(_0307_ ), .B2(_0594_ ), .ZN(_0623_ ) );
OAI21_X1 _1316_ ( .A(_0534_ ), .B1(_0622_ ), .B2(_0623_ ), .ZN(_0624_ ) );
NAND3_X1 _1317_ ( .A1(_0375_ ), .A2(_0602_ ), .A3(_0292_ ), .ZN(_0625_ ) );
AOI21_X1 _1318_ ( .A(_0533_ ), .B1(_0624_ ), .B2(_0625_ ), .ZN(_0626_ ) );
OAI22_X1 _1319_ ( .A1(_0583_ ), .A2(_0278_ ), .B1(_0335_ ), .B2(_0594_ ), .ZN(_0627_ ) );
OAI21_X1 _1320_ ( .A(_0300_ ), .B1(_0626_ ), .B2(_0627_ ), .ZN(_0628_ ) );
NAND3_X1 _1321_ ( .A1(_0375_ ), .A2(_0602_ ), .A3(_0277_ ), .ZN(_0629_ ) );
AOI21_X1 _1322_ ( .A(_0285_ ), .B1(_0628_ ), .B2(_0629_ ), .ZN(_0630_ ) );
OAI21_X1 _1323_ ( .A(_0259_ ), .B1(_0560_ ), .B2(_0352_ ), .ZN(_0631_ ) );
OAI211_X1 _1324_ ( .A(_0631_ ), .B(_0331_ ), .C1(_0278_ ), .C2(_0594_ ), .ZN(_0632_ ) );
OAI21_X1 _1325_ ( .A(_0532_ ), .B1(_0630_ ), .B2(_0632_ ), .ZN(_0633_ ) );
NAND3_X1 _1326_ ( .A1(_0375_ ), .A2(_0602_ ), .A3(_0259_ ), .ZN(_0634_ ) );
AOI21_X1 _1327_ ( .A(_0512_ ), .B1(_0633_ ), .B2(_0634_ ), .ZN(_0635_ ) );
NAND3_X1 _1328_ ( .A1(_0375_ ), .A2(_0602_ ), .A3(_0325_ ), .ZN(_0636_ ) );
AND3_X1 _1329_ ( .A1(_0369_ ), .A2(_0351_ ), .A3(_0259_ ), .ZN(_0637_ ) );
AOI21_X1 _1330_ ( .A(_0389_ ), .B1(_0364_ ), .B2(_0308_ ), .ZN(_0638_ ) );
AOI211_X1 _1331_ ( .A(_0637_ ), .B(_0638_ ), .C1(_0325_ ), .C2(_0582_ ), .ZN(_0639_ ) );
OAI21_X1 _1332_ ( .A(_0636_ ), .B1(_0639_ ), .B2(_0387_ ), .ZN(_0640_ ) );
OAI21_X1 _1333_ ( .A(_0514_ ), .B1(_0635_ ), .B2(_0640_ ), .ZN(_0641_ ) );
AND3_X1 _1334_ ( .A1(_0369_ ), .A2(_0351_ ), .A3(_0325_ ), .ZN(_0642_ ) );
INV_X1 _1335_ ( .A(_0642_ ), .ZN(_0643_ ) );
AOI21_X1 _1336_ ( .A(reset ), .B1(_0641_ ), .B2(_0643_ ), .ZN(_0042_ ) );
NAND2_X1 _1337_ ( .A1(_0314_ ), .A2(_0362_ ), .ZN(_0644_ ) );
OAI21_X1 _1338_ ( .A(_0444_ ), .B1(_0644_ ), .B2(_0355_ ), .ZN(_0645_ ) );
AND2_X1 _1339_ ( .A1(_0645_ ), .A2(_0482_ ), .ZN(_0646_ ) );
AOI21_X1 _1340_ ( .A(_0492_ ), .B1(_0471_ ), .B2(_0404_ ), .ZN(_0647_ ) );
AND2_X1 _1341_ ( .A1(_0273_ ), .A2(_0404_ ), .ZN(_0648_ ) );
AOI221_X4 _1342_ ( .A(_0648_ ), .B1(_0302_ ), .B2(_0397_ ), .C1(_0333_ ), .C2(_0404_ ), .ZN(_0649_ ) );
OAI211_X1 _1343_ ( .A(_0375_ ), .B(_0371_ ), .C1(_0397_ ), .C2(_0399_ ), .ZN(_0650_ ) );
NAND2_X1 _1344_ ( .A1(_0644_ ), .A2(_0385_ ), .ZN(_0651_ ) );
AND4_X1 _1345_ ( .A1(_0647_ ), .A2(_0649_ ), .A3(_0650_ ), .A4(_0651_ ), .ZN(_0652_ ) );
AOI211_X1 _1346_ ( .A(\inst_o[7] ), .B(_0317_ ), .C1(_0274_ ), .C2(_0362_ ), .ZN(_0653_ ) );
AOI211_X1 _1347_ ( .A(_0496_ ), .B(_0653_ ), .C1(_0471_ ), .C2(_0467_ ), .ZN(_0654_ ) );
OAI21_X1 _1348_ ( .A(_0644_ ), .B1(_0438_ ), .B2(_0495_ ), .ZN(_0655_ ) );
AND4_X1 _1349_ ( .A1(_0646_ ), .A2(_0652_ ), .A3(_0654_ ), .A4(_0655_ ), .ZN(_0656_ ) );
AOI21_X1 _1350_ ( .A(_0386_ ), .B1(_0471_ ), .B2(_0399_ ), .ZN(_0657_ ) );
NOR3_X1 _1351_ ( .A1(_0332_ ), .A2(_0271_ ), .A3(_0638_ ), .ZN(_0658_ ) );
OAI21_X1 _1352_ ( .A(_0516_ ), .B1(_0644_ ), .B2(_0355_ ), .ZN(_0659_ ) );
OAI21_X1 _1353_ ( .A(_0265_ ), .B1(_0644_ ), .B2(_0355_ ), .ZN(_0660_ ) );
AND4_X1 _1354_ ( .A1(_0657_ ), .A2(_0658_ ), .A3(_0659_ ), .A4(_0660_ ), .ZN(_0661_ ) );
AOI211_X1 _1355_ ( .A(reset ), .B(_0642_ ), .C1(_0656_ ), .C2(_0661_ ), .ZN(_0043_ ) );
OAI21_X1 _1356_ ( .A(_0580_ ), .B1(_0049_ ), .B2(_0317_ ), .ZN(_0662_ ) );
NOR4_X1 _1357_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0663_ ) );
NAND4_X1 _1358_ ( .A1(_0663_ ), .A2(_0210_ ), .A3(_0214_ ), .A4(_0215_ ), .ZN(_0664_ ) );
NOR2_X1 _1359_ ( .A1(_0664_ ), .A2(_0047_ ), .ZN(_0665_ ) );
AND4_X1 _1360_ ( .A1(_0316_ ), .A2(_0053_ ), .A3(\i5.io_mem_data[3] ), .A4(_0291_ ), .ZN(_0666_ ) );
OAI211_X1 _1361_ ( .A(_0662_ ), .B(_0665_ ), .C1(\i0.io_Pc_count[3] ), .C2(_0666_ ), .ZN(_0667_ ) );
NAND2_X1 _1362_ ( .A1(_0662_ ), .A2(_0226_ ), .ZN(_0668_ ) );
NOR4_X1 _1363_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0669_ ) );
NOR4_X1 _1364_ ( .A1(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0670_ ) );
NOR4_X1 _1365_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0671_ ) );
NOR4_X1 _1366_ ( .A1(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .A4(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0672_ ) );
NAND4_X1 _1367_ ( .A1(_0669_ ), .A2(_0670_ ), .A3(_0671_ ), .A4(_0672_ ), .ZN(_0673_ ) );
INV_X1 _1368_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_0674_ ) );
NAND4_X1 _1369_ ( .A1(_0674_ ), .A2(\i0.io_Pc_count[15] ), .A3(\inst_o[2] ), .A4(\inst_o[0] ), .ZN(_0675_ ) );
OR3_X1 _1370_ ( .A1(_0673_ ), .A2(_0202_ ), .A3(_0675_ ), .ZN(_0676_ ) );
NOR4_X1 _1371_ ( .A1(_0667_ ), .A2(_0668_ ), .A3(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .A4(_0676_ ), .ZN(ALU_carry ) );
NOR2_X1 _1372_ ( .A1(_0667_ ), .A2(_0676_ ), .ZN(_0677_ ) );
AND4_X1 _1373_ ( .A1(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .A2(_0677_ ), .A3(_0226_ ), .A4(_0662_ ), .ZN(ALU_overflow ) );
AOI221_X4 _1374_ ( .A(_0125_ ), .B1(_0053_ ), .B2(_0385_ ), .C1(\inst_o[3] ), .C2(_0243_ ), .ZN(\i0.state_$_SDFFE_PP0P__Q_E ) );
AOI22_X1 _1375_ ( .A1(_0243_ ), .A2(\inst_o[3] ), .B1(_0053_ ), .B2(_0385_ ), .ZN(\i0.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
CLKGATE_X1 _1376_ ( .CK(clk ), .E(\i0.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_0678_ ) );
CLKGATE_X1 _1377_ ( .CK(clk ), .E(\i0.state_$_SDFFE_PP0P__Q_E ), .GCK(_0679_ ) );
LOGIC0_X1 _1378_ ( .Z(\inst_o[10] ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q ( .D(_0000_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[10] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_1 ( .D(_0001_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[9] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_10 ( .D(_0002_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[29] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_11 ( .D(_0003_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[28] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_12 ( .D(_0004_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[27] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_13 ( .D(_0005_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[26] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_14 ( .D(_0006_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[25] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_15 ( .D(_0007_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[24] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_16 ( .D(_0008_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[23] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_17 ( .D(_0009_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[22] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_18 ( .D(_0010_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[21] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_19 ( .D(_0011_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[20] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_2 ( .D(_0012_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[8] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_20 ( .D(_0013_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[19] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_21 ( .D(_0014_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[18] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_22 ( .D(_0015_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[17] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_23 ( .D(_0016_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[16] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_24 ( .D(_0017_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[15] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_25 ( .D(_0018_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[14] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_26 ( .D(_0019_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[13] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_27 ( .D(_0020_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[12] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_28 ( .D(_0021_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[11] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_3 ( .D(_0022_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[7] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_4 ( .D(_0023_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[6] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_5 ( .D(_0024_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[5] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_6 ( .D(_0025_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[4] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_7 ( .D(_0026_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[3] ), .QN(_0693_ ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_8 ( .D(_0027_ ), .CK(_0679_ ), .Q(\i0.io_Pc_count[2] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_9 ( .D(_0028_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[30] ), .QN(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP1P__Q ( .D(_0029_ ), .CK(_0678_ ), .Q(\i0.io_Pc_count[31] ), .QN(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q ( .D(_0030_ ), .CK(clk ), .Q(\inst_o[7] ), .QN(_0692_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_1 ( .D(_0031_ ), .CK(clk ), .Q(\inst_o[6] ), .QN(_0691_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_2 ( .D(_0032_ ), .CK(clk ), .Q(\inst_o[5] ), .QN(_0690_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_3 ( .D(_0033_ ), .CK(clk ), .Q(\inst_o[4] ), .QN(_0689_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_4 ( .D(_0034_ ), .CK(clk ), .Q(\inst_o[3] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XNOR__A_Y_$_NAND__A_B ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_5 ( .D(_0035_ ), .CK(clk ), .Q(\inst_o[2] ), .QN(_0688_ ) );
DFF_X1 \i1.data1_$_SDFF_PP0__Q_6 ( .D(\inst_o[10] ), .CK(clk ), .Q(\inst_o[0] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_ORNOT__Y_A_$_ORNOT__Y_B_$_XOR__A_Y_$_OR__A_1_B ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q ( .D(_0036_ ), .CK(clk ), .Q(\i5.io_mem_data[7] ), .QN(_0687_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_1 ( .D(_0037_ ), .CK(clk ), .Q(\i5.io_mem_data[6] ), .QN(_0686_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_2 ( .D(_0038_ ), .CK(clk ), .Q(\i5.io_mem_data[5] ), .QN(_0685_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_3 ( .D(_0039_ ), .CK(clk ), .Q(\i5.io_mem_data[4] ), .QN(_0684_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_4 ( .D(_0040_ ), .CK(clk ), .Q(\i5.io_mem_data[3] ), .QN(_0683_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_5 ( .D(_0041_ ), .CK(clk ), .Q(\i5.io_mem_data[2] ), .QN(_0682_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_6 ( .D(_0042_ ), .CK(clk ), .Q(\i5.io_mem_data[1] ), .QN(_0681_ ) );
DFF_X1 \i9.data1_$_SDFF_PP0__Q_7 ( .D(_0043_ ), .CK(clk ), .Q(\i5.io_mem_data[0] ), .QN(_0680_ ) );

endmodule
