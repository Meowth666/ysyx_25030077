module MyOperators(
  input         clock,
  input         reset,
  input  [31:0] io_instruction,
  input  [31:0] io_rs1_data,
  input  [31:0] io_rs2_data,
  input  [31:0] io_imm_data,
  output [31:0] io_mem_data
);
  wire [7:0] _index_T_2 = io_instruction[7:0] ^ io_rs1_data[7:0]; // @[module.scala 15:35]
  wire [7:0] _index_T_4 = _index_T_2 ^ io_rs2_data[7:0]; // @[module.scala 15:54]
  wire [7:0] index = _index_T_4 ^ io_imm_data[7:0]; // @[module.scala 15:73]
  wire [31:0] _GEN_1 = 8'h1 == index ? 32'h1 : 32'h0; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_2 = 8'h2 == index ? 32'h2 : _GEN_1; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_3 = 8'h3 == index ? 32'h3 : _GEN_2; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_4 = 8'h4 == index ? 32'h4 : _GEN_3; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_5 = 8'h5 == index ? 32'h5 : _GEN_4; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_6 = 8'h6 == index ? 32'h6 : _GEN_5; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_7 = 8'h7 == index ? 32'h7 : _GEN_6; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_8 = 8'h8 == index ? 32'h8 : _GEN_7; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_9 = 8'h9 == index ? 32'h9 : _GEN_8; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_10 = 8'ha == index ? 32'ha : _GEN_9; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_11 = 8'hb == index ? 32'hb : _GEN_10; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_12 = 8'hc == index ? 32'hc : _GEN_11; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_13 = 8'hd == index ? 32'hd : _GEN_12; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_14 = 8'he == index ? 32'he : _GEN_13; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_15 = 8'hf == index ? 32'hf : _GEN_14; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_16 = 8'h10 == index ? 32'h10 : _GEN_15; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_17 = 8'h11 == index ? 32'h11 : _GEN_16; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_18 = 8'h12 == index ? 32'h12 : _GEN_17; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_19 = 8'h13 == index ? 32'h13 : _GEN_18; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_20 = 8'h14 == index ? 32'h14 : _GEN_19; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_21 = 8'h15 == index ? 32'h15 : _GEN_20; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_22 = 8'h16 == index ? 32'h16 : _GEN_21; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_23 = 8'h17 == index ? 32'h17 : _GEN_22; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_24 = 8'h18 == index ? 32'h18 : _GEN_23; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_25 = 8'h19 == index ? 32'h19 : _GEN_24; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_26 = 8'h1a == index ? 32'h1a : _GEN_25; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_27 = 8'h1b == index ? 32'h1b : _GEN_26; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_28 = 8'h1c == index ? 32'h1c : _GEN_27; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_29 = 8'h1d == index ? 32'h1d : _GEN_28; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_30 = 8'h1e == index ? 32'h1e : _GEN_29; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_31 = 8'h1f == index ? 32'h1f : _GEN_30; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_32 = 8'h20 == index ? 32'h20 : _GEN_31; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_33 = 8'h21 == index ? 32'h21 : _GEN_32; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_34 = 8'h22 == index ? 32'h22 : _GEN_33; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_35 = 8'h23 == index ? 32'h23 : _GEN_34; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_36 = 8'h24 == index ? 32'h24 : _GEN_35; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_37 = 8'h25 == index ? 32'h25 : _GEN_36; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_38 = 8'h26 == index ? 32'h26 : _GEN_37; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_39 = 8'h27 == index ? 32'h27 : _GEN_38; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_40 = 8'h28 == index ? 32'h28 : _GEN_39; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_41 = 8'h29 == index ? 32'h29 : _GEN_40; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_42 = 8'h2a == index ? 32'h2a : _GEN_41; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_43 = 8'h2b == index ? 32'h2b : _GEN_42; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_44 = 8'h2c == index ? 32'h2c : _GEN_43; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_45 = 8'h2d == index ? 32'h2d : _GEN_44; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_46 = 8'h2e == index ? 32'h2e : _GEN_45; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_47 = 8'h2f == index ? 32'h2f : _GEN_46; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_48 = 8'h30 == index ? 32'h30 : _GEN_47; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_49 = 8'h31 == index ? 32'h31 : _GEN_48; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_50 = 8'h32 == index ? 32'h32 : _GEN_49; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_51 = 8'h33 == index ? 32'h33 : _GEN_50; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_52 = 8'h34 == index ? 32'h34 : _GEN_51; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_53 = 8'h35 == index ? 32'h35 : _GEN_52; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_54 = 8'h36 == index ? 32'h36 : _GEN_53; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_55 = 8'h37 == index ? 32'h37 : _GEN_54; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_56 = 8'h38 == index ? 32'h38 : _GEN_55; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_57 = 8'h39 == index ? 32'h39 : _GEN_56; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_58 = 8'h3a == index ? 32'h3a : _GEN_57; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_59 = 8'h3b == index ? 32'h3b : _GEN_58; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_60 = 8'h3c == index ? 32'h3c : _GEN_59; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_61 = 8'h3d == index ? 32'h3d : _GEN_60; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_62 = 8'h3e == index ? 32'h3e : _GEN_61; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_63 = 8'h3f == index ? 32'h3f : _GEN_62; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_64 = 8'h40 == index ? 32'h40 : _GEN_63; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_65 = 8'h41 == index ? 32'h41 : _GEN_64; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_66 = 8'h42 == index ? 32'h42 : _GEN_65; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_67 = 8'h43 == index ? 32'h43 : _GEN_66; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_68 = 8'h44 == index ? 32'h44 : _GEN_67; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_69 = 8'h45 == index ? 32'h45 : _GEN_68; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_70 = 8'h46 == index ? 32'h46 : _GEN_69; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_71 = 8'h47 == index ? 32'h47 : _GEN_70; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_72 = 8'h48 == index ? 32'h48 : _GEN_71; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_73 = 8'h49 == index ? 32'h49 : _GEN_72; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_74 = 8'h4a == index ? 32'h4a : _GEN_73; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_75 = 8'h4b == index ? 32'h4b : _GEN_74; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_76 = 8'h4c == index ? 32'h4c : _GEN_75; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_77 = 8'h4d == index ? 32'h4d : _GEN_76; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_78 = 8'h4e == index ? 32'h4e : _GEN_77; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_79 = 8'h4f == index ? 32'h4f : _GEN_78; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_80 = 8'h50 == index ? 32'h50 : _GEN_79; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_81 = 8'h51 == index ? 32'h51 : _GEN_80; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_82 = 8'h52 == index ? 32'h52 : _GEN_81; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_83 = 8'h53 == index ? 32'h53 : _GEN_82; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_84 = 8'h54 == index ? 32'h54 : _GEN_83; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_85 = 8'h55 == index ? 32'h55 : _GEN_84; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_86 = 8'h56 == index ? 32'h56 : _GEN_85; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_87 = 8'h57 == index ? 32'h57 : _GEN_86; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_88 = 8'h58 == index ? 32'h58 : _GEN_87; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_89 = 8'h59 == index ? 32'h59 : _GEN_88; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_90 = 8'h5a == index ? 32'h5a : _GEN_89; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_91 = 8'h5b == index ? 32'h5b : _GEN_90; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_92 = 8'h5c == index ? 32'h5c : _GEN_91; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_93 = 8'h5d == index ? 32'h5d : _GEN_92; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_94 = 8'h5e == index ? 32'h5e : _GEN_93; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_95 = 8'h5f == index ? 32'h5f : _GEN_94; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_96 = 8'h60 == index ? 32'h60 : _GEN_95; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_97 = 8'h61 == index ? 32'h61 : _GEN_96; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_98 = 8'h62 == index ? 32'h62 : _GEN_97; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_99 = 8'h63 == index ? 32'h63 : _GEN_98; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_100 = 8'h64 == index ? 32'h64 : _GEN_99; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_101 = 8'h65 == index ? 32'h65 : _GEN_100; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_102 = 8'h66 == index ? 32'h66 : _GEN_101; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_103 = 8'h67 == index ? 32'h67 : _GEN_102; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_104 = 8'h68 == index ? 32'h68 : _GEN_103; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_105 = 8'h69 == index ? 32'h69 : _GEN_104; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_106 = 8'h6a == index ? 32'h6a : _GEN_105; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_107 = 8'h6b == index ? 32'h6b : _GEN_106; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_108 = 8'h6c == index ? 32'h6c : _GEN_107; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_109 = 8'h6d == index ? 32'h6d : _GEN_108; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_110 = 8'h6e == index ? 32'h6e : _GEN_109; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_111 = 8'h6f == index ? 32'h6f : _GEN_110; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_112 = 8'h70 == index ? 32'h70 : _GEN_111; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_113 = 8'h71 == index ? 32'h71 : _GEN_112; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_114 = 8'h72 == index ? 32'h72 : _GEN_113; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_115 = 8'h73 == index ? 32'h73 : _GEN_114; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_116 = 8'h74 == index ? 32'h74 : _GEN_115; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_117 = 8'h75 == index ? 32'h75 : _GEN_116; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_118 = 8'h76 == index ? 32'h76 : _GEN_117; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_119 = 8'h77 == index ? 32'h77 : _GEN_118; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_120 = 8'h78 == index ? 32'h78 : _GEN_119; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_121 = 8'h79 == index ? 32'h79 : _GEN_120; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_122 = 8'h7a == index ? 32'h7a : _GEN_121; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_123 = 8'h7b == index ? 32'h7b : _GEN_122; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_124 = 8'h7c == index ? 32'h7c : _GEN_123; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_125 = 8'h7d == index ? 32'h7d : _GEN_124; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_126 = 8'h7e == index ? 32'h7e : _GEN_125; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_127 = 8'h7f == index ? 32'h7f : _GEN_126; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_128 = 8'h80 == index ? 32'h80 : _GEN_127; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_129 = 8'h81 == index ? 32'h81 : _GEN_128; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_130 = 8'h82 == index ? 32'h82 : _GEN_129; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_131 = 8'h83 == index ? 32'h83 : _GEN_130; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_132 = 8'h84 == index ? 32'h84 : _GEN_131; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_133 = 8'h85 == index ? 32'h85 : _GEN_132; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_134 = 8'h86 == index ? 32'h86 : _GEN_133; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_135 = 8'h87 == index ? 32'h87 : _GEN_134; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_136 = 8'h88 == index ? 32'h88 : _GEN_135; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_137 = 8'h89 == index ? 32'h89 : _GEN_136; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_138 = 8'h8a == index ? 32'h8a : _GEN_137; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_139 = 8'h8b == index ? 32'h8b : _GEN_138; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_140 = 8'h8c == index ? 32'h8c : _GEN_139; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_141 = 8'h8d == index ? 32'h8d : _GEN_140; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_142 = 8'h8e == index ? 32'h8e : _GEN_141; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_143 = 8'h8f == index ? 32'h8f : _GEN_142; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_144 = 8'h90 == index ? 32'h90 : _GEN_143; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_145 = 8'h91 == index ? 32'h91 : _GEN_144; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_146 = 8'h92 == index ? 32'h92 : _GEN_145; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_147 = 8'h93 == index ? 32'h93 : _GEN_146; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_148 = 8'h94 == index ? 32'h94 : _GEN_147; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_149 = 8'h95 == index ? 32'h95 : _GEN_148; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_150 = 8'h96 == index ? 32'h96 : _GEN_149; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_151 = 8'h97 == index ? 32'h97 : _GEN_150; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_152 = 8'h98 == index ? 32'h98 : _GEN_151; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_153 = 8'h99 == index ? 32'h99 : _GEN_152; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_154 = 8'h9a == index ? 32'h9a : _GEN_153; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_155 = 8'h9b == index ? 32'h9b : _GEN_154; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_156 = 8'h9c == index ? 32'h9c : _GEN_155; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_157 = 8'h9d == index ? 32'h9d : _GEN_156; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_158 = 8'h9e == index ? 32'h9e : _GEN_157; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_159 = 8'h9f == index ? 32'h9f : _GEN_158; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_160 = 8'ha0 == index ? 32'ha0 : _GEN_159; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_161 = 8'ha1 == index ? 32'ha1 : _GEN_160; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_162 = 8'ha2 == index ? 32'ha2 : _GEN_161; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_163 = 8'ha3 == index ? 32'ha3 : _GEN_162; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_164 = 8'ha4 == index ? 32'ha4 : _GEN_163; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_165 = 8'ha5 == index ? 32'ha5 : _GEN_164; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_166 = 8'ha6 == index ? 32'ha6 : _GEN_165; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_167 = 8'ha7 == index ? 32'ha7 : _GEN_166; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_168 = 8'ha8 == index ? 32'ha8 : _GEN_167; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_169 = 8'ha9 == index ? 32'ha9 : _GEN_168; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_170 = 8'haa == index ? 32'haa : _GEN_169; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_171 = 8'hab == index ? 32'hab : _GEN_170; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_172 = 8'hac == index ? 32'hac : _GEN_171; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_173 = 8'had == index ? 32'had : _GEN_172; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_174 = 8'hae == index ? 32'hae : _GEN_173; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_175 = 8'haf == index ? 32'haf : _GEN_174; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_176 = 8'hb0 == index ? 32'hb0 : _GEN_175; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_177 = 8'hb1 == index ? 32'hb1 : _GEN_176; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_178 = 8'hb2 == index ? 32'hb2 : _GEN_177; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_179 = 8'hb3 == index ? 32'hb3 : _GEN_178; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_180 = 8'hb4 == index ? 32'hb4 : _GEN_179; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_181 = 8'hb5 == index ? 32'hb5 : _GEN_180; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_182 = 8'hb6 == index ? 32'hb6 : _GEN_181; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_183 = 8'hb7 == index ? 32'hb7 : _GEN_182; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_184 = 8'hb8 == index ? 32'hb8 : _GEN_183; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_185 = 8'hb9 == index ? 32'hb9 : _GEN_184; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_186 = 8'hba == index ? 32'hba : _GEN_185; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_187 = 8'hbb == index ? 32'hbb : _GEN_186; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_188 = 8'hbc == index ? 32'hbc : _GEN_187; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_189 = 8'hbd == index ? 32'hbd : _GEN_188; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_190 = 8'hbe == index ? 32'hbe : _GEN_189; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_191 = 8'hbf == index ? 32'hbf : _GEN_190; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_192 = 8'hc0 == index ? 32'hc0 : _GEN_191; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_193 = 8'hc1 == index ? 32'hc1 : _GEN_192; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_194 = 8'hc2 == index ? 32'hc2 : _GEN_193; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_195 = 8'hc3 == index ? 32'hc3 : _GEN_194; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_196 = 8'hc4 == index ? 32'hc4 : _GEN_195; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_197 = 8'hc5 == index ? 32'hc5 : _GEN_196; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_198 = 8'hc6 == index ? 32'hc6 : _GEN_197; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_199 = 8'hc7 == index ? 32'hc7 : _GEN_198; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_200 = 8'hc8 == index ? 32'hc8 : _GEN_199; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_201 = 8'hc9 == index ? 32'hc9 : _GEN_200; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_202 = 8'hca == index ? 32'hca : _GEN_201; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_203 = 8'hcb == index ? 32'hcb : _GEN_202; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_204 = 8'hcc == index ? 32'hcc : _GEN_203; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_205 = 8'hcd == index ? 32'hcd : _GEN_204; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_206 = 8'hce == index ? 32'hce : _GEN_205; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_207 = 8'hcf == index ? 32'hcf : _GEN_206; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_208 = 8'hd0 == index ? 32'hd0 : _GEN_207; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_209 = 8'hd1 == index ? 32'hd1 : _GEN_208; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_210 = 8'hd2 == index ? 32'hd2 : _GEN_209; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_211 = 8'hd3 == index ? 32'hd3 : _GEN_210; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_212 = 8'hd4 == index ? 32'hd4 : _GEN_211; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_213 = 8'hd5 == index ? 32'hd5 : _GEN_212; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_214 = 8'hd6 == index ? 32'hd6 : _GEN_213; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_215 = 8'hd7 == index ? 32'hd7 : _GEN_214; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_216 = 8'hd8 == index ? 32'hd8 : _GEN_215; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_217 = 8'hd9 == index ? 32'hd9 : _GEN_216; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_218 = 8'hda == index ? 32'hda : _GEN_217; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_219 = 8'hdb == index ? 32'hdb : _GEN_218; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_220 = 8'hdc == index ? 32'hdc : _GEN_219; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_221 = 8'hdd == index ? 32'hdd : _GEN_220; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_222 = 8'hde == index ? 32'hde : _GEN_221; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_223 = 8'hdf == index ? 32'hdf : _GEN_222; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_224 = 8'he0 == index ? 32'he0 : _GEN_223; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_225 = 8'he1 == index ? 32'he1 : _GEN_224; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_226 = 8'he2 == index ? 32'he2 : _GEN_225; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_227 = 8'he3 == index ? 32'he3 : _GEN_226; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_228 = 8'he4 == index ? 32'he4 : _GEN_227; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_229 = 8'he5 == index ? 32'he5 : _GEN_228; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_230 = 8'he6 == index ? 32'he6 : _GEN_229; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_231 = 8'he7 == index ? 32'he7 : _GEN_230; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_232 = 8'he8 == index ? 32'he8 : _GEN_231; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_233 = 8'he9 == index ? 32'he9 : _GEN_232; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_234 = 8'hea == index ? 32'hea : _GEN_233; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_235 = 8'heb == index ? 32'heb : _GEN_234; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_236 = 8'hec == index ? 32'hec : _GEN_235; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_237 = 8'hed == index ? 32'hed : _GEN_236; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_238 = 8'hee == index ? 32'hee : _GEN_237; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_239 = 8'hef == index ? 32'hef : _GEN_238; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_240 = 8'hf0 == index ? 32'hf0 : _GEN_239; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_241 = 8'hf1 == index ? 32'hf1 : _GEN_240; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_242 = 8'hf2 == index ? 32'hf2 : _GEN_241; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_243 = 8'hf3 == index ? 32'hf3 : _GEN_242; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_244 = 8'hf4 == index ? 32'hf4 : _GEN_243; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_245 = 8'hf5 == index ? 32'hf5 : _GEN_244; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_246 = 8'hf6 == index ? 32'hf6 : _GEN_245; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_247 = 8'hf7 == index ? 32'hf7 : _GEN_246; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_248 = 8'hf8 == index ? 32'hf8 : _GEN_247; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_249 = 8'hf9 == index ? 32'hf9 : _GEN_248; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_250 = 8'hfa == index ? 32'hfa : _GEN_249; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_251 = 8'hfb == index ? 32'hfb : _GEN_250; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_252 = 8'hfc == index ? 32'hfc : _GEN_251; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_253 = 8'hfd == index ? 32'hfd : _GEN_252; // @[module.scala 17:{15,15}]
  wire [31:0] _GEN_254 = 8'hfe == index ? 32'hfe : _GEN_253; // @[module.scala 17:{15,15}]
  assign io_mem_data = 8'hff == index ? 32'hff : _GEN_254; // @[module.scala 17:{15,15}]
endmodule
