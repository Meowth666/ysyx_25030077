//Generate the verilog at 2025-08-31T15:58:11 by iSTA.
module ysyx_25030077_top (
clk,
reset,
ALU_carry,
ALU_overflow,
PC_count_o
);

input clk ;
input reset ;
output ALU_carry ;
output ALU_overflow ;
output [31:0] PC_count_o ;

wire clk ;
wire reset ;
wire ALU_carry ;
wire ALU_overflow ;
wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_AND__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XOR__A_B_$_OR__B_Y_$_OR__B_Y_$_NOR__A_B_$_ORNOT__A_Y_$_ORNOT__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_NAND__B_1_Y_$_ORNOT__A_Y_$_ANDNOT__A_1_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ;
wire ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_A_$_OR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \PC_count_o[0] ;
wire \PC_count_o[1] ;
wire \PC_count_o[2] ;
wire \PC_count_o[3] ;
wire \PC_count_o[4] ;
wire \PC_count_o[5] ;
wire \PC_count_o[6] ;
wire \PC_count_o[7] ;
wire \PC_count_o[8] ;
wire \PC_count_o[9] ;
wire \PC_count_o[10] ;
wire \PC_count_o[11] ;
wire \PC_count_o[12] ;
wire \PC_count_o[13] ;
wire \PC_count_o[14] ;
wire \PC_count_o[15] ;
wire \PC_count_o[16] ;
wire \PC_count_o[17] ;
wire \PC_count_o[18] ;
wire \PC_count_o[19] ;
wire \PC_count_o[20] ;
wire \PC_count_o[21] ;
wire \PC_count_o[22] ;
wire \PC_count_o[23] ;
wire \PC_count_o[24] ;
wire \PC_count_o[25] ;
wire \PC_count_o[26] ;
wire \PC_count_o[27] ;
wire \PC_count_o[28] ;
wire \PC_count_o[29] ;
wire \PC_count_o[30] ;
wire \PC_count_o[31] ;

assign ALU_carry = ALU_overflow ;
assign ALU_carry = \PC_count_o[0] ;
assign ALU_carry = \PC_count_o[1] ;
assign PC_count_o[2] = \PC_count_o[2] ;
assign PC_count_o[3] = \PC_count_o[3] ;
assign PC_count_o[4] = \PC_count_o[4] ;
assign PC_count_o[5] = \PC_count_o[5] ;
assign PC_count_o[6] = \PC_count_o[6] ;
assign PC_count_o[7] = \PC_count_o[7] ;
assign PC_count_o[8] = \PC_count_o[8] ;
assign PC_count_o[9] = \PC_count_o[9] ;
assign PC_count_o[10] = \PC_count_o[10] ;
assign PC_count_o[11] = \PC_count_o[11] ;
assign PC_count_o[12] = \PC_count_o[12] ;
assign PC_count_o[13] = \PC_count_o[13] ;
assign PC_count_o[14] = \PC_count_o[14] ;
assign PC_count_o[15] = \PC_count_o[15] ;
assign PC_count_o[16] = \PC_count_o[16] ;
assign PC_count_o[17] = \PC_count_o[17] ;
assign PC_count_o[18] = \PC_count_o[18] ;
assign PC_count_o[19] = \PC_count_o[19] ;
assign PC_count_o[20] = \PC_count_o[20] ;
assign PC_count_o[21] = \PC_count_o[21] ;
assign PC_count_o[22] = \PC_count_o[22] ;
assign PC_count_o[23] = \PC_count_o[23] ;
assign PC_count_o[24] = \PC_count_o[24] ;
assign PC_count_o[25] = \PC_count_o[25] ;
assign PC_count_o[26] = \PC_count_o[26] ;
assign PC_count_o[27] = \PC_count_o[27] ;
assign PC_count_o[28] = \PC_count_o[28] ;
assign PC_count_o[29] = \PC_count_o[29] ;
assign PC_count_o[30] = \PC_count_o[30] ;
assign PC_count_o[31] = \PC_count_o[31] ;

AND2_X4 _135_ ( .A1(\PC_count_o[3] ), .A2(\PC_count_o[2] ), .ZN(_126_ ) );
AND2_X4 _136_ ( .A1(\PC_count_o[5] ), .A2(\PC_count_o[4] ), .ZN(_127_ ) );
AND2_X4 _137_ ( .A1(_126_ ), .A2(_127_ ), .ZN(_128_ ) );
AND4_X1 _138_ ( .A1(\PC_count_o[7] ), .A2(\PC_count_o[6] ), .A3(\PC_count_o[9] ), .A4(\PC_count_o[8] ), .ZN(_129_ ) );
AND2_X4 _139_ ( .A1(_128_ ), .A2(_129_ ), .ZN(_130_ ) );
INV_X1 _140_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_131_ ) );
AND2_X1 _141_ ( .A1(_130_ ), .A2(_131_ ), .ZN(_030_ ) );
INV_X1 _142_ ( .A(reset ), .ZN(_031_ ) );
OAI21_X1 _143_ ( .A(_031_ ), .B1(_130_ ), .B2(_131_ ), .ZN(_032_ ) );
NOR2_X1 _144_ ( .A1(_030_ ), .A2(_032_ ), .ZN(_000_ ) );
NAND3_X1 _145_ ( .A1(_128_ ), .A2(\PC_count_o[7] ), .A3(\PC_count_o[6] ), .ZN(_033_ ) );
NOR2_X1 _146_ ( .A1(_033_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_034_ ) );
XNOR2_X1 _147_ ( .A(_034_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_035_ ) );
CLKBUF_X2 _148_ ( .A(_031_ ), .Z(_036_ ) );
AND2_X1 _149_ ( .A1(_035_ ), .A2(_036_ ), .ZN(_001_ ) );
AND2_X4 _150_ ( .A1(\PC_count_o[13] ), .A2(\PC_count_o[12] ), .ZN(_037_ ) );
AND3_X4 _151_ ( .A1(_037_ ), .A2(\PC_count_o[11] ), .A3(\PC_count_o[10] ), .ZN(_038_ ) );
AND2_X1 _152_ ( .A1(\PC_count_o[15] ), .A2(\PC_count_o[14] ), .ZN(_039_ ) );
AND4_X4 _153_ ( .A1(\PC_count_o[16] ), .A2(_038_ ), .A3(\PC_count_o[17] ), .A4(_039_ ), .ZN(_040_ ) );
AND2_X4 _154_ ( .A1(_040_ ), .A2(_130_ ), .ZN(_041_ ) );
AND4_X1 _155_ ( .A1(\PC_count_o[24] ), .A2(\PC_count_o[23] ), .A3(\PC_count_o[25] ), .A4(\PC_count_o[22] ), .ZN(_042_ ) );
AND2_X1 _156_ ( .A1(\PC_count_o[19] ), .A2(\PC_count_o[18] ), .ZN(_043_ ) );
AND4_X1 _157_ ( .A1(\PC_count_o[20] ), .A2(_042_ ), .A3(\PC_count_o[21] ), .A4(_043_ ), .ZN(_044_ ) );
AND2_X4 _158_ ( .A1(_041_ ), .A2(_044_ ), .ZN(_045_ ) );
NAND3_X4 _159_ ( .A1(_045_ ), .A2(\PC_count_o[27] ), .A3(\PC_count_o[26] ), .ZN(_046_ ) );
OR3_X4 _160_ ( .A1(_046_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_047_ ) );
OAI21_X1 _161_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_046_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_048_ ) );
AND3_X1 _162_ ( .A1(_047_ ), .A2(_036_ ), .A3(_048_ ), .ZN(_002_ ) );
NOR2_X1 _163_ ( .A1(_046_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_049_ ) );
INV_X1 _164_ ( .A(_049_ ), .ZN(_050_ ) );
AOI21_X1 _165_ ( .A(reset ), .B1(_046_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_051_ ) );
AND2_X1 _166_ ( .A1(_050_ ), .A2(_051_ ), .ZN(_003_ ) );
INV_X1 _167_ ( .A(_045_ ), .ZN(_052_ ) );
OR3_X4 _168_ ( .A1(_052_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_053_ ) );
OAI21_X1 _169_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_052_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_054_ ) );
AND3_X1 _170_ ( .A1(_053_ ), .A2(_036_ ), .A3(_054_ ), .ZN(_004_ ) );
NOR2_X1 _171_ ( .A1(_052_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_055_ ) );
INV_X1 _172_ ( .A(_055_ ), .ZN(_056_ ) );
AOI21_X1 _173_ ( .A(reset ), .B1(_052_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_057_ ) );
AND2_X1 _174_ ( .A1(_056_ ), .A2(_057_ ), .ZN(_005_ ) );
AND3_X1 _175_ ( .A1(_043_ ), .A2(\PC_count_o[20] ), .A3(\PC_count_o[21] ), .ZN(_058_ ) );
AND3_X4 _176_ ( .A1(_040_ ), .A2(_130_ ), .A3(_058_ ), .ZN(_059_ ) );
AND3_X4 _177_ ( .A1(_059_ ), .A2(\PC_count_o[23] ), .A3(\PC_count_o[22] ), .ZN(_060_ ) );
INV_X2 _178_ ( .A(_060_ ), .ZN(_061_ ) );
OR3_X4 _179_ ( .A1(_061_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_062_ ) );
OAI21_X1 _180_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_061_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_063_ ) );
AND3_X1 _181_ ( .A1(_062_ ), .A2(_036_ ), .A3(_063_ ), .ZN(_006_ ) );
NOR2_X1 _182_ ( .A1(_061_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_064_ ) );
INV_X1 _183_ ( .A(_064_ ), .ZN(_065_ ) );
AOI21_X1 _184_ ( .A(reset ), .B1(_061_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_066_ ) );
AND2_X1 _185_ ( .A1(_065_ ), .A2(_066_ ), .ZN(_007_ ) );
INV_X1 _186_ ( .A(_059_ ), .ZN(_067_ ) );
OR3_X1 _187_ ( .A1(_067_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_068_ ) );
OAI21_X1 _188_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_067_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_069_ ) );
AND3_X1 _189_ ( .A1(_068_ ), .A2(_036_ ), .A3(_069_ ), .ZN(_008_ ) );
NOR2_X1 _190_ ( .A1(_067_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_070_ ) );
INV_X1 _191_ ( .A(_070_ ), .ZN(_071_ ) );
AOI21_X1 _192_ ( .A(reset ), .B1(_067_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_072_ ) );
AND2_X1 _193_ ( .A1(_071_ ), .A2(_072_ ), .ZN(_009_ ) );
NAND3_X1 _194_ ( .A1(_040_ ), .A2(_130_ ), .A3(_043_ ), .ZN(_073_ ) );
OR3_X1 _195_ ( .A1(_073_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_074_ ) );
OAI21_X1 _196_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_073_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_075_ ) );
AND3_X1 _197_ ( .A1(_074_ ), .A2(_036_ ), .A3(_075_ ), .ZN(_010_ ) );
NOR2_X1 _198_ ( .A1(_073_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_076_ ) );
INV_X1 _199_ ( .A(_076_ ), .ZN(_077_ ) );
AOI21_X1 _200_ ( .A(reset ), .B1(_073_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_078_ ) );
AND2_X1 _201_ ( .A1(_077_ ), .A2(_078_ ), .ZN(_011_ ) );
INV_X1 _202_ ( .A(_034_ ), .ZN(_079_ ) );
AOI21_X1 _203_ ( .A(reset ), .B1(_033_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_080_ ) );
AND2_X1 _204_ ( .A1(_079_ ), .A2(_080_ ), .ZN(_012_ ) );
INV_X1 _205_ ( .A(_041_ ), .ZN(_081_ ) );
OR3_X1 _206_ ( .A1(_081_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_082_ ) );
OAI21_X1 _207_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_081_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_083_ ) );
AND3_X1 _208_ ( .A1(_082_ ), .A2(_036_ ), .A3(_083_ ), .ZN(_013_ ) );
NOR2_X1 _209_ ( .A1(_081_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_084_ ) );
INV_X1 _210_ ( .A(_084_ ), .ZN(_085_ ) );
AOI21_X1 _211_ ( .A(reset ), .B1(_081_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_086_ ) );
AND2_X1 _212_ ( .A1(_085_ ), .A2(_086_ ), .ZN(_014_ ) );
AND3_X1 _213_ ( .A1(_130_ ), .A2(_038_ ), .A3(_039_ ), .ZN(_087_ ) );
INV_X1 _214_ ( .A(_087_ ), .ZN(_088_ ) );
OR3_X1 _215_ ( .A1(_088_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_089_ ) );
OAI21_X1 _216_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_088_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_090_ ) );
AND3_X1 _217_ ( .A1(_089_ ), .A2(_036_ ), .A3(_090_ ), .ZN(_015_ ) );
AND3_X1 _218_ ( .A1(_130_ ), .A2(\PC_count_o[11] ), .A3(\PC_count_o[10] ), .ZN(_091_ ) );
NAND3_X1 _219_ ( .A1(_091_ ), .A2(_037_ ), .A3(_039_ ), .ZN(_092_ ) );
OR2_X1 _220_ ( .A1(_092_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_093_ ) );
AOI21_X1 _221_ ( .A(reset ), .B1(_088_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_094_ ) );
AND2_X1 _222_ ( .A1(_093_ ), .A2(_094_ ), .ZN(_016_ ) );
AND3_X1 _223_ ( .A1(_038_ ), .A2(_128_ ), .A3(_129_ ), .ZN(_095_ ) );
INV_X1 _224_ ( .A(_095_ ), .ZN(_096_ ) );
OR3_X1 _225_ ( .A1(_096_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_097_ ) );
OAI21_X1 _226_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_096_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_098_ ) );
AND3_X1 _227_ ( .A1(_097_ ), .A2(_031_ ), .A3(_098_ ), .ZN(_017_ ) );
NAND2_X1 _228_ ( .A1(_091_ ), .A2(_037_ ), .ZN(_099_ ) );
OR2_X1 _229_ ( .A1(_099_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_100_ ) );
AOI21_X1 _230_ ( .A(reset ), .B1(_096_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_101_ ) );
AND2_X1 _231_ ( .A1(_100_ ), .A2(_101_ ), .ZN(_018_ ) );
INV_X1 _232_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_102_ ) );
AND2_X1 _233_ ( .A1(_091_ ), .A2(_102_ ), .ZN(_103_ ) );
OR2_X1 _234_ ( .A1(_103_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_104_ ) );
NAND3_X1 _235_ ( .A1(_091_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(_102_ ), .ZN(_105_ ) );
AOI21_X1 _236_ ( .A(reset ), .B1(_104_ ), .B2(_105_ ), .ZN(_019_ ) );
OAI21_X1 _237_ ( .A(_031_ ), .B1(_091_ ), .B2(_102_ ), .ZN(_106_ ) );
NOR2_X1 _238_ ( .A1(_103_ ), .A2(_106_ ), .ZN(_020_ ) );
INV_X1 _239_ ( .A(_030_ ), .ZN(_107_ ) );
AOI21_X1 _240_ ( .A(reset ), .B1(_107_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_A_$_OR__Y_B ), .ZN(_108_ ) );
INV_X1 _241_ ( .A(_130_ ), .ZN(_109_ ) );
OR3_X1 _242_ ( .A1(_109_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_A_$_OR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_110_ ) );
AND2_X1 _243_ ( .A1(_108_ ), .A2(_110_ ), .ZN(_021_ ) );
INV_X1 _244_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_111_ ) );
AND2_X1 _245_ ( .A1(_128_ ), .A2(_111_ ), .ZN(_112_ ) );
XNOR2_X1 _246_ ( .A(_112_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_113_ ) );
AND2_X1 _247_ ( .A1(_113_ ), .A2(_036_ ), .ZN(_022_ ) );
OAI21_X1 _248_ ( .A(_031_ ), .B1(_128_ ), .B2(_111_ ), .ZN(_114_ ) );
NOR2_X1 _249_ ( .A1(_112_ ), .A2(_114_ ), .ZN(_023_ ) );
INV_X1 _250_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_115_ ) );
AND2_X1 _251_ ( .A1(_126_ ), .A2(_115_ ), .ZN(_116_ ) );
XNOR2_X1 _252_ ( .A(_116_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_117_ ) );
AND2_X1 _253_ ( .A1(_117_ ), .A2(_036_ ), .ZN(_024_ ) );
OAI21_X1 _254_ ( .A(_031_ ), .B1(_126_ ), .B2(_115_ ), .ZN(_118_ ) );
NOR2_X1 _255_ ( .A1(_116_ ), .A2(_118_ ), .ZN(_025_ ) );
NOR2_X1 _256_ ( .A1(\PC_count_o[3] ), .A2(\PC_count_o[2] ), .ZN(_119_ ) );
NOR3_X1 _257_ ( .A1(_126_ ), .A2(_119_ ), .A3(reset ), .ZN(_026_ ) );
NOR2_X1 _258_ ( .A1(reset ), .A2(\PC_count_o[2] ), .ZN(_027_ ) );
AND4_X1 _259_ ( .A1(\PC_count_o[29] ), .A2(\PC_count_o[28] ), .A3(\PC_count_o[27] ), .A4(\PC_count_o[26] ), .ZN(_120_ ) );
NAND3_X1 _260_ ( .A1(_041_ ), .A2(_044_ ), .A3(_120_ ), .ZN(_121_ ) );
NOR2_X1 _261_ ( .A1(_121_ ), .A2(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_122_ ) );
INV_X1 _262_ ( .A(_122_ ), .ZN(_123_ ) );
AOI21_X1 _263_ ( .A(reset ), .B1(_121_ ), .B2(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_124_ ) );
AND2_X1 _264_ ( .A1(_123_ ), .A2(_124_ ), .ZN(_028_ ) );
AOI21_X1 _265_ ( .A(reset ), .B1(_122_ ), .B2(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_125_ ) );
OAI21_X1 _266_ ( .A(_125_ ), .B1(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_122_ ), .ZN(_029_ ) );
CLKGATE_X1 _267_ ( .CK(clk ), .E(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_AND__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XOR__A_B_$_OR__B_Y_$_OR__B_Y_$_NOR__A_B_$_ORNOT__A_Y_$_ORNOT__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_NAND__B_1_Y_$_ORNOT__A_Y_$_ANDNOT__A_1_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_132_ ) );
CLKGATE_X1 _268_ ( .CK(clk ), .E(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_AND__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XOR__A_B_$_OR__B_Y_$_OR__B_Y_$_NOR__A_B_$_ORNOT__A_Y_$_ORNOT__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_NAND__B_1_Y_$_ORNOT__A_Y_$_ANDNOT__A_1_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_133_ ) );
LOGIC1_X1 _269_ ( .Z(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_A_$_AND__Y_B_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_XOR__A_B_$_OR__B_Y_$_OR__B_Y_$_NOR__A_B_$_ORNOT__A_Y_$_ORNOT__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_NAND__B_1_Y_$_ORNOT__A_Y_$_ANDNOT__A_1_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
LOGIC0_X1 _270_ ( .Z(ALU_carry ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q ( .D(_000_ ), .CK(_133_ ), .Q(\PC_count_o[10] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_1 ( .D(_001_ ), .CK(_133_ ), .Q(\PC_count_o[9] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_10 ( .D(_002_ ), .CK(_132_ ), .Q(\PC_count_o[29] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_11 ( .D(_003_ ), .CK(_132_ ), .Q(\PC_count_o[28] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_12 ( .D(_004_ ), .CK(_132_ ), .Q(\PC_count_o[27] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_13 ( .D(_005_ ), .CK(_132_ ), .Q(\PC_count_o[26] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_14 ( .D(_006_ ), .CK(_132_ ), .Q(\PC_count_o[25] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_15 ( .D(_007_ ), .CK(_132_ ), .Q(\PC_count_o[24] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_16 ( .D(_008_ ), .CK(_132_ ), .Q(\PC_count_o[23] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_17 ( .D(_009_ ), .CK(_132_ ), .Q(\PC_count_o[22] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_18 ( .D(_010_ ), .CK(_132_ ), .Q(\PC_count_o[21] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_19 ( .D(_011_ ), .CK(_132_ ), .Q(\PC_count_o[20] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_2 ( .D(_012_ ), .CK(_133_ ), .Q(\PC_count_o[8] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_20 ( .D(_013_ ), .CK(_132_ ), .Q(\PC_count_o[19] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_21 ( .D(_014_ ), .CK(_132_ ), .Q(\PC_count_o[18] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_22 ( .D(_015_ ), .CK(_132_ ), .Q(\PC_count_o[17] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_23 ( .D(_016_ ), .CK(_132_ ), .Q(\PC_count_o[16] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_24 ( .D(_017_ ), .CK(_132_ ), .Q(\PC_count_o[15] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_25 ( .D(_018_ ), .CK(_132_ ), .Q(\PC_count_o[14] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_26 ( .D(_019_ ), .CK(_132_ ), .Q(\PC_count_o[13] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_27 ( .D(_020_ ), .CK(_132_ ), .Q(\PC_count_o[12] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_28 ( .D(_021_ ), .CK(_132_ ), .Q(\PC_count_o[11] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_B_$_XOR__Y_A_$_OR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_3 ( .D(_022_ ), .CK(_133_ ), .Q(\PC_count_o[7] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_4 ( .D(_023_ ), .CK(_133_ ), .Q(\PC_count_o[6] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_5 ( .D(_024_ ), .CK(_133_ ), .Q(\PC_count_o[5] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_6 ( .D(_025_ ), .CK(_133_ ), .Q(\PC_count_o[4] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_7 ( .D(_026_ ), .CK(_133_ ), .Q(\PC_count_o[3] ), .QN(_134_ ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_8 ( .D(_027_ ), .CK(_133_ ), .Q(\PC_count_o[2] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_9 ( .D(_028_ ), .CK(_132_ ), .Q(\PC_count_o[30] ), .QN(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP1P__Q ( .D(_029_ ), .CK(_132_ ), .Q(\PC_count_o[31] ), .QN(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ) );

endmodule
