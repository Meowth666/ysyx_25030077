module ysyx_25030077_IDU(
  input  [31:0] io_instruction,
  output [2:0]  io_imm_type,
  output [4:0]  io_rs1,
  output [4:0]  io_rs2,
  output [4:0]  io_rd,
  output [2:0]  io_data_control,
  output [3:0]  io_ALU_ctrl,
  output [3:0]  io_pc_next_type,
  output [2:0]  io_r_mask,
  output [2:0]  io_w_mask,
  output        io_r_valid,        
  output        is_break_out
);

  assign is_break_out = (io_instruction == 32'h100073);
  
  wire [4:0] addi_Rs1 = io_instruction[19:15]; // @[IDU.scala 30:32]
  wire [4:0] addi_Rd = io_instruction[11:7]; // @[IDU.scala 31:32]
  wire [4:0] sltu_Rs2 = io_instruction[24:20]; // @[IDU.scala 96:33]
  wire [9:0] _isaddi_T_2 = {io_instruction[14:12],io_instruction[6:0]}; // @[Cat.scala 31:58]
  wire  isaddi = _isaddi_T_2 == 10'h13; // @[IDU.scala 294:64]
  wire  isxori = _isaddi_T_2 == 10'h213; // @[IDU.scala 295:64]
  wire  isori = _isaddi_T_2 == 10'h313; // @[IDU.scala 296:64]
  wire  isandi = _isaddi_T_2 == 10'h393; // @[IDU.scala 297:64]
  wire [15:0] _issrai_T_3 = {io_instruction[31:26],io_instruction[14:12],io_instruction[6:0]}; // @[Cat.scala 31:58]
  wire  issrai = _issrai_T_3 == 16'h4293; // @[IDU.scala 298:87]
  wire  issrli = _issrai_T_3 == 16'h293; // @[IDU.scala 299:87]
  wire  isslli = _issrai_T_3 == 16'h93; // @[IDU.scala 300:87]
  wire  issra = _issrai_T_3 == 16'h42b3; // @[IDU.scala 301:87]
  wire  issrl = _issrai_T_3 == 16'h2b3; // @[IDU.scala 302:87]
  wire  isbeq = _isaddi_T_2 == 10'h63; // @[IDU.scala 303:64]
  wire  isbne = _isaddi_T_2 == 10'he3; // @[IDU.scala 304:64]
  wire [16:0] _isadd_T_3 = {io_instruction[31:25],io_instruction[14:12],io_instruction[6:0]}; // @[Cat.scala 31:58]
  wire  isadd = _isadd_T_3 == 17'h33; // @[IDU.scala 305:87]
  wire  isxor = _isadd_T_3 == 17'h233; // @[IDU.scala 306:87]
  wire  isand = _isadd_T_3 == 17'h3b3; // @[IDU.scala 307:87]
  wire  isor = _isadd_T_3 == 17'h333; // @[IDU.scala 308:87]
  wire  issub = _isadd_T_3 == 17'h8033; // @[IDU.scala 309:87]
  wire  islui = io_instruction[6:0] == 7'h37; // @[IDU.scala 310:36]
  wire  isauipc = io_instruction[6:0] == 7'h17; // @[IDU.scala 311:38]
  wire  isjal = io_instruction[6:0] == 7'h6f; // @[IDU.scala 312:36]
  wire  isjalr = _isaddi_T_2 == 10'h67; // @[IDU.scala 313:65]
  wire  issw = _isaddi_T_2 == 10'h123; // @[IDU.scala 314:63]
  wire  isbge = _isaddi_T_2 == 10'h2e3; // @[IDU.scala 315:63]
  wire  isblt = _isaddi_T_2 == 10'h263; // @[IDU.scala 316:63]
  wire  isbltu = _isaddi_T_2 == 10'h363; // @[IDU.scala 317:63]
  wire  isbgeu = _isaddi_T_2 == 10'h3e3; // @[IDU.scala 318:63]
  wire  issb = _isaddi_T_2 == 10'h23; // @[IDU.scala 319:63]
  wire  issh = _isaddi_T_2 == 10'ha3; // @[IDU.scala 320:63]
  wire  islbu = _isaddi_T_2 == 10'h203; // @[IDU.scala 321:63]
  wire  islb = _isaddi_T_2 == 10'h3; // @[IDU.scala 322:63]
  wire  islw = _isaddi_T_2 == 10'h103; // @[IDU.scala 323:63]
  wire  islh = _isaddi_T_2 == 10'h83; // @[IDU.scala 324:63]
  wire  islhu = _isaddi_T_2 == 10'h283; // @[IDU.scala 325:63]
  wire  issll = _isadd_T_3 == 17'hb3; // @[IDU.scala 326:86]
  wire  isslt = _isadd_T_3 == 17'h133; // @[IDU.scala 327:88]
  wire  issltu = _isadd_T_3 == 17'h1b3; // @[IDU.scala 328:88]
  wire  issltiu = _isaddi_T_2 == 10'h193; // @[IDU.scala 329:65]
  wire  isslti = _isaddi_T_2 == 10'h113; // @[IDU.scala 330:65]
  wire  iscsrrw = _isaddi_T_2 == 10'hf3; // @[IDU.scala 331:67]
  wire  iscsrrs = _isaddi_T_2 == 10'h173; // @[IDU.scala 332:67]
  wire  isebreak = io_instruction == 32'h100073; // @[IDU.scala 333:34]
  wire  isecall = io_instruction == 32'h73; // @[IDU.scala 334:34]
  wire  ismret = io_instruction == 32'h30200073; // @[IDU.scala 335:34]
  wire [2:0] _io_imm_type_T = islb ? 3'h1 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_1 = islbu ? 3'h1 : _io_imm_type_T; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_2 = islhu ? 3'h1 : _io_imm_type_T_1; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_3 = islh ? 3'h1 : _io_imm_type_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_4 = islw ? 3'h1 : _io_imm_type_T_3; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_5 = issh ? 3'h4 : _io_imm_type_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_6 = issb ? 3'h4 : _io_imm_type_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_7 = issw ? 3'h4 : _io_imm_type_T_6; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_8 = isjalr ? 3'h3 : _io_imm_type_T_7; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_9 = isjal ? 3'h3 : _io_imm_type_T_8; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_10 = isauipc ? 3'h2 : _io_imm_type_T_9; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_11 = islui ? 3'h2 : _io_imm_type_T_10; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_12 = isslti ? 3'h1 : _io_imm_type_T_11; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_13 = issltiu ? 3'h1 : _io_imm_type_T_12; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_14 = isslli ? 3'h5 : _io_imm_type_T_13; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_15 = issrli ? 3'h5 : _io_imm_type_T_14; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_16 = issrai ? 3'h5 : _io_imm_type_T_15; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_17 = iscsrrs ? 3'h6 : _io_imm_type_T_16; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_18 = iscsrrw ? 3'h6 : _io_imm_type_T_17; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_19 = isandi ? 3'h1 : _io_imm_type_T_18; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_20 = isori ? 3'h1 : _io_imm_type_T_19; // @[Mux.scala 101:16]
  wire [2:0] _io_imm_type_T_21 = isxori ? 3'h1 : _io_imm_type_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T = isslt ? addi_Rs1 : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_1 = issltu ? addi_Rs1 : _io_rs1_T; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_2 = isbne ? addi_Rs1 : _io_rs1_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_3 = isbgeu ? addi_Rs1 : _io_rs1_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_4 = isbltu ? addi_Rs1 : _io_rs1_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_5 = isblt ? addi_Rs1 : _io_rs1_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_6 = isbge ? addi_Rs1 : _io_rs1_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_7 = isbeq ? addi_Rs1 : _io_rs1_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_8 = issub ? addi_Rs1 : _io_rs1_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_9 = isor ? addi_Rs1 : _io_rs1_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_10 = isxor ? addi_Rs1 : _io_rs1_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_11 = issrl ? addi_Rs1 : _io_rs1_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_12 = issra ? addi_Rs1 : _io_rs1_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_13 = issll ? addi_Rs1 : _io_rs1_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_14 = isand ? addi_Rs1 : _io_rs1_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_15 = isadd ? addi_Rs1 : _io_rs1_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_16 = islb ? addi_Rs1 : _io_rs1_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_17 = islbu ? addi_Rs1 : _io_rs1_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_18 = islhu ? addi_Rs1 : _io_rs1_T_17; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_19 = islh ? addi_Rs1 : _io_rs1_T_18; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_20 = islw ? addi_Rs1 : _io_rs1_T_19; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_21 = issh ? addi_Rs1 : _io_rs1_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_22 = issb ? addi_Rs1 : _io_rs1_T_21; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_23 = issw ? addi_Rs1 : _io_rs1_T_22; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_24 = isjalr ? addi_Rs1 : _io_rs1_T_23; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_25 = isslti ? addi_Rs1 : _io_rs1_T_24; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_26 = issltiu ? addi_Rs1 : _io_rs1_T_25; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_27 = isslli ? addi_Rs1 : _io_rs1_T_26; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_28 = issrli ? addi_Rs1 : _io_rs1_T_27; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_29 = issrai ? addi_Rs1 : _io_rs1_T_28; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_30 = iscsrrs ? addi_Rs1 : _io_rs1_T_29; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_31 = iscsrrw ? addi_Rs1 : _io_rs1_T_30; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_32 = isandi ? addi_Rs1 : _io_rs1_T_31; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_33 = isori ? addi_Rs1 : _io_rs1_T_32; // @[Mux.scala 101:16]
  wire [4:0] _io_rs1_T_34 = isxori ? addi_Rs1 : _io_rs1_T_33; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T = isslt ? sltu_Rs2 : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_1 = issltu ? sltu_Rs2 : _io_rs2_T; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_2 = isbne ? sltu_Rs2 : _io_rs2_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_3 = isbgeu ? sltu_Rs2 : _io_rs2_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_4 = isbltu ? sltu_Rs2 : _io_rs2_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_5 = isblt ? sltu_Rs2 : _io_rs2_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_6 = isbge ? sltu_Rs2 : _io_rs2_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_7 = isbeq ? sltu_Rs2 : _io_rs2_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_8 = issub ? sltu_Rs2 : _io_rs2_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_9 = isor ? sltu_Rs2 : _io_rs2_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_10 = isxor ? sltu_Rs2 : _io_rs2_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_11 = issrl ? sltu_Rs2 : _io_rs2_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_12 = issra ? sltu_Rs2 : _io_rs2_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_13 = issll ? sltu_Rs2 : _io_rs2_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_14 = isand ? sltu_Rs2 : _io_rs2_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_15 = isadd ? sltu_Rs2 : _io_rs2_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_16 = issh ? sltu_Rs2 : _io_rs2_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_rs2_T_17 = issb ? sltu_Rs2 : _io_rs2_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T = isslt ? addi_Rd : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_1 = issltu ? addi_Rd : _io_rd_T; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_2 = issub ? addi_Rd : _io_rd_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_3 = isor ? addi_Rd : _io_rd_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_4 = isxor ? addi_Rd : _io_rd_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_5 = issrl ? addi_Rd : _io_rd_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_6 = issra ? addi_Rd : _io_rd_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_7 = issll ? addi_Rd : _io_rd_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_8 = isand ? addi_Rd : _io_rd_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_9 = isadd ? addi_Rd : _io_rd_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_10 = islb ? addi_Rd : _io_rd_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_11 = islbu ? addi_Rd : _io_rd_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_12 = islhu ? addi_Rd : _io_rd_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_13 = islh ? addi_Rd : _io_rd_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_14 = islw ? addi_Rd : _io_rd_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_15 = isjalr ? addi_Rd : _io_rd_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_16 = isjal ? addi_Rd : _io_rd_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_17 = isauipc ? addi_Rd : _io_rd_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_18 = islui ? addi_Rd : _io_rd_T_17; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_19 = isslti ? addi_Rd : _io_rd_T_18; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_20 = issltiu ? addi_Rd : _io_rd_T_19; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_21 = isslli ? addi_Rd : _io_rd_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_22 = issrli ? addi_Rd : _io_rd_T_21; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_23 = issrai ? addi_Rd : _io_rd_T_22; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_24 = iscsrrs ? addi_Rd : _io_rd_T_23; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_25 = iscsrrw ? addi_Rd : _io_rd_T_24; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_26 = isandi ? addi_Rd : _io_rd_T_25; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_27 = isori ? addi_Rd : _io_rd_T_26; // @[Mux.scala 101:16]
  wire [4:0] _io_rd_T_28 = isxori ? addi_Rd : _io_rd_T_27; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T = issltu ? 5'h2 : 5'h0; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_1 = isslt ? 5'ha : _io_ALU_ctrl_T; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_2 = isbne ? 5'h0 : _io_ALU_ctrl_T_1; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_3 = isbgeu ? 5'h0 : _io_ALU_ctrl_T_2; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_4 = isbltu ? 5'h0 : _io_ALU_ctrl_T_3; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_5 = isblt ? 5'h0 : _io_ALU_ctrl_T_4; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_6 = isbge ? 5'h0 : _io_ALU_ctrl_T_5; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_7 = isbeq ? 5'h0 : _io_ALU_ctrl_T_6; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_8 = issub ? 5'h1 : _io_ALU_ctrl_T_7; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_9 = isor ? 5'h3 : _io_ALU_ctrl_T_8; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_10 = isxor ? 5'h4 : _io_ALU_ctrl_T_9; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_11 = issrl ? 5'h9 : _io_ALU_ctrl_T_10; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_12 = issra ? 5'h5 : _io_ALU_ctrl_T_11; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_13 = issll ? 5'h8 : _io_ALU_ctrl_T_12; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_14 = isand ? 5'h6 : _io_ALU_ctrl_T_13; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_15 = isadd ? 5'h0 : _io_ALU_ctrl_T_14; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_16 = islb ? 5'h0 : _io_ALU_ctrl_T_15; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_17 = islbu ? 5'h0 : _io_ALU_ctrl_T_16; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_18 = islhu ? 5'h0 : _io_ALU_ctrl_T_17; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_19 = islh ? 5'h0 : _io_ALU_ctrl_T_18; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_20 = islw ? 5'h0 : _io_ALU_ctrl_T_19; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_21 = issh ? 5'h0 : _io_ALU_ctrl_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_22 = issb ? 5'h0 : _io_ALU_ctrl_T_21; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_23 = issw ? 5'h0 : _io_ALU_ctrl_T_22; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_24 = isjalr ? 5'h0 : _io_ALU_ctrl_T_23; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_25 = isjal ? 5'h0 : _io_ALU_ctrl_T_24; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_26 = isauipc ? 5'h0 : _io_ALU_ctrl_T_25; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_27 = islui ? 5'h0 : _io_ALU_ctrl_T_26; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_28 = isslti ? 5'ha : _io_ALU_ctrl_T_27; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_29 = issltiu ? 5'h2 : _io_ALU_ctrl_T_28; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_30 = isslli ? 5'h8 : _io_ALU_ctrl_T_29; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_31 = issrli ? 5'h9 : _io_ALU_ctrl_T_30; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_32 = issrai ? 5'h5 : _io_ALU_ctrl_T_31; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_33 = iscsrrs ? 5'hc : _io_ALU_ctrl_T_32; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_34 = iscsrrw ? 5'hb : _io_ALU_ctrl_T_33; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_35 = isandi ? 5'h6 : _io_ALU_ctrl_T_34; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_36 = isori ? 5'h3 : _io_ALU_ctrl_T_35; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_37 = isxori ? 5'h4 : _io_ALU_ctrl_T_36; // @[Mux.scala 101:16]
  wire [4:0] _io_ALU_ctrl_T_38 = isaddi ? 5'h0 : _io_ALU_ctrl_T_37; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T = issltu ? 3'h3 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_1 = isslt ? 3'h3 : _io_data_control_T; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_2 = isbne ? 3'h0 : _io_data_control_T_1; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_3 = isbgeu ? 3'h0 : _io_data_control_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_4 = isbltu ? 3'h0 : _io_data_control_T_3; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_5 = isblt ? 3'h0 : _io_data_control_T_4; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_6 = isbge ? 3'h0 : _io_data_control_T_5; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_7 = isbeq ? 3'h0 : _io_data_control_T_6; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_8 = issub ? 3'h3 : _io_data_control_T_7; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_9 = isor ? 3'h3 : _io_data_control_T_8; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_10 = isxor ? 3'h3 : _io_data_control_T_9; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_11 = issrl ? 3'h3 : _io_data_control_T_10; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_12 = issra ? 3'h3 : _io_data_control_T_11; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_13 = issll ? 3'h3 : _io_data_control_T_12; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_14 = isand ? 3'h3 : _io_data_control_T_13; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_15 = isadd ? 3'h3 : _io_data_control_T_14; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_16 = islb ? 3'h2 : _io_data_control_T_15; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_17 = islbu ? 3'h2 : _io_data_control_T_16; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_18 = islhu ? 3'h2 : _io_data_control_T_17; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_19 = islh ? 3'h2 : _io_data_control_T_18; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_20 = islw ? 3'h2 : _io_data_control_T_19; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_21 = issh ? 3'h0 : _io_data_control_T_20; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_22 = issb ? 3'h0 : _io_data_control_T_21; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_23 = issw ? 3'h0 : _io_data_control_T_22; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_24 = isjalr ? 3'h1 : _io_data_control_T_23; // @[Mux.scala 101:16]
  wire [2:0] _io_data_control_T_25 = isjal ? 3'h1 : _io_data_control_T_24; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T = isslti ? 4'h0 : 4'h3; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_1 = issltiu ? 4'h0 : _io_pc_next_type_T; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_2 = isslt ? 4'h0 : _io_pc_next_type_T_1; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_3 = issltu ? 4'h0 : _io_pc_next_type_T_2; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_4 = isbne ? 4'h5 : _io_pc_next_type_T_3; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_5 = isbgeu ? 4'h8 : _io_pc_next_type_T_4; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_6 = isbltu ? 4'ha : _io_pc_next_type_T_5; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_7 = isblt ? 4'h9 : _io_pc_next_type_T_6; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_8 = isbge ? 4'h7 : _io_pc_next_type_T_7; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_9 = isbeq ? 4'h6 : _io_pc_next_type_T_8; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_10 = issub ? 4'h0 : _io_pc_next_type_T_9; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_11 = isor ? 4'h0 : _io_pc_next_type_T_10; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_12 = isxor ? 4'h0 : _io_pc_next_type_T_11; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_13 = issrl ? 4'h0 : _io_pc_next_type_T_12; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_14 = issra ? 4'h0 : _io_pc_next_type_T_13; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_15 = issll ? 4'h0 : _io_pc_next_type_T_14; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_16 = isand ? 4'h0 : _io_pc_next_type_T_15; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_17 = isadd ? 4'h0 : _io_pc_next_type_T_16; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_18 = islb ? 4'h0 : _io_pc_next_type_T_17; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_19 = islbu ? 4'h0 : _io_pc_next_type_T_18; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_20 = islhu ? 4'h0 : _io_pc_next_type_T_19; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_21 = islh ? 4'h0 : _io_pc_next_type_T_20; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_22 = islw ? 4'h0 : _io_pc_next_type_T_21; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_23 = ismret ? 4'hc : _io_pc_next_type_T_22; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_24 = isecall ? 4'hb : _io_pc_next_type_T_23; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_25 = isebreak ? 4'h4 : _io_pc_next_type_T_24; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_26 = issh ? 4'h0 : _io_pc_next_type_T_25; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_27 = issb ? 4'h0 : _io_pc_next_type_T_26; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_28 = issw ? 4'h0 : _io_pc_next_type_T_27; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_29 = isslli ? 4'h0 : _io_pc_next_type_T_28; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_30 = issrli ? 4'h0 : _io_pc_next_type_T_29; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_31 = issrai ? 4'h0 : _io_pc_next_type_T_30; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_32 = iscsrrs ? 4'h0 : _io_pc_next_type_T_31; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_33 = iscsrrw ? 4'h0 : _io_pc_next_type_T_32; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_34 = isandi ? 4'h0 : _io_pc_next_type_T_33; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_35 = isori ? 4'h0 : _io_pc_next_type_T_34; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_36 = isxori ? 4'h0 : _io_pc_next_type_T_35; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_37 = isaddi ? 4'h0 : _io_pc_next_type_T_36; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_38 = islui ? 4'h0 : _io_pc_next_type_T_37; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_39 = isauipc ? 4'h0 : _io_pc_next_type_T_38; // @[Mux.scala 101:16]
  wire [3:0] _io_pc_next_type_T_40 = isjalr ? 4'h2 : _io_pc_next_type_T_39; // @[Mux.scala 101:16]
  wire [2:0] _io_r_mask_T = islb ? 3'h5 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_r_mask_T_1 = islbu ? 3'h2 : _io_r_mask_T; // @[Mux.scala 101:16]
  wire [2:0] _io_r_mask_T_2 = islhu ? 3'h4 : _io_r_mask_T_1; // @[Mux.scala 101:16]
  wire [2:0] _io_r_mask_T_3 = islh ? 3'h3 : _io_r_mask_T_2; // @[Mux.scala 101:16]
  wire [2:0] _io_w_mask_T = issh ? 3'h2 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _io_w_mask_T_1 = issb ? 3'h3 : _io_w_mask_T; // @[Mux.scala 101:16]
  assign io_imm_type = isaddi ? 3'h1 : _io_imm_type_T_21; // @[Mux.scala 101:16]
  assign io_rs1 = isaddi ? addi_Rs1 : _io_rs1_T_34; // @[Mux.scala 101:16]
  assign io_rs2 = issw ? sltu_Rs2 : _io_rs2_T_17; // @[Mux.scala 101:16]
  assign io_rd = isaddi ? addi_Rd : _io_rd_T_28; // @[Mux.scala 101:16]
  assign io_data_control = isauipc ? 3'h1 : _io_data_control_T_25; // @[Mux.scala 101:16]
  assign io_ALU_ctrl = _io_ALU_ctrl_T_38[3:0]; // @[IDU.scala 458:15]
  assign io_pc_next_type = isjal ? 4'h1 : _io_pc_next_type_T_40; // @[Mux.scala 101:16]
  assign io_r_mask = islw ? 3'h1 : _io_r_mask_T_3; // @[Mux.scala 101:16]
  assign io_w_mask = issw ? 3'h1 : _io_w_mask_T_1; // @[Mux.scala 101:16]
  assign io_r_valid = islw | (islh | (islhu | (islbu | islb))); // @[Mux.scala 101:16]
endmodule
