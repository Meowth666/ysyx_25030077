//Generate the verilog at 2025-08-31T15:22:19 by iSTA.
module ysyx_25030077_top (
clk,
reset,
ALU_carry,
ALU_overflow,
imm,
rd,
ALU_ctrl,
rs1_out,
rs2_out,
PC_count_o
);

input clk ;
input reset ;
output ALU_carry ;
output ALU_overflow ;
output [31:0] imm ;
output [4:0] rd ;
output [3:0] ALU_ctrl ;
output [31:0] rs1_out ;
output [31:0] rs2_out ;
output [31:0] PC_count_o ;

wire clk ;
wire reset ;
wire ALU_carry ;
wire ALU_overflow ;
wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ;
wire ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ;
wire \i0.state_$_SDFFE_PP0P__Q_E ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ;
wire \imm[0] ;
wire \imm[1] ;
wire \imm[2] ;
wire \imm[3] ;
wire \imm[4] ;
wire \imm[5] ;
wire \imm[6] ;
wire \imm[7] ;
wire \imm[8] ;
wire \imm[9] ;
wire \imm[10] ;
wire \imm[11] ;
wire \imm[12] ;
wire \imm[13] ;
wire \imm[14] ;
wire \imm[15] ;
wire \imm[16] ;
wire \imm[17] ;
wire \imm[18] ;
wire \imm[19] ;
wire \imm[20] ;
wire \imm[21] ;
wire \imm[22] ;
wire \imm[23] ;
wire \imm[24] ;
wire \imm[25] ;
wire \imm[26] ;
wire \imm[27] ;
wire \imm[28] ;
wire \imm[29] ;
wire \imm[30] ;
wire \imm[31] ;
wire \rd[0] ;
wire \rd[1] ;
wire \rd[2] ;
wire \rd[3] ;
wire \rd[4] ;
wire \ALU_ctrl[0] ;
wire \ALU_ctrl[1] ;
wire \ALU_ctrl[2] ;
wire \ALU_ctrl[3] ;
wire \rs1_out[0] ;
wire \rs1_out[1] ;
wire \rs1_out[2] ;
wire \rs1_out[3] ;
wire \rs1_out[4] ;
wire \rs1_out[5] ;
wire \rs1_out[6] ;
wire \rs1_out[7] ;
wire \rs1_out[8] ;
wire \rs1_out[9] ;
wire \rs1_out[10] ;
wire \rs1_out[11] ;
wire \rs1_out[12] ;
wire \rs1_out[13] ;
wire \rs1_out[14] ;
wire \rs1_out[15] ;
wire \rs1_out[16] ;
wire \rs1_out[17] ;
wire \rs1_out[18] ;
wire \rs1_out[19] ;
wire \rs1_out[20] ;
wire \rs1_out[21] ;
wire \rs1_out[22] ;
wire \rs1_out[23] ;
wire \rs1_out[24] ;
wire \rs1_out[25] ;
wire \rs1_out[26] ;
wire \rs1_out[27] ;
wire \rs1_out[28] ;
wire \rs1_out[29] ;
wire \rs1_out[30] ;
wire \rs1_out[31] ;
wire \rs2_out[0] ;
wire \rs2_out[1] ;
wire \rs2_out[2] ;
wire \rs2_out[3] ;
wire \rs2_out[4] ;
wire \rs2_out[5] ;
wire \rs2_out[6] ;
wire \rs2_out[7] ;
wire \rs2_out[8] ;
wire \rs2_out[9] ;
wire \rs2_out[10] ;
wire \rs2_out[11] ;
wire \rs2_out[12] ;
wire \rs2_out[13] ;
wire \rs2_out[14] ;
wire \rs2_out[15] ;
wire \rs2_out[16] ;
wire \rs2_out[17] ;
wire \rs2_out[18] ;
wire \rs2_out[19] ;
wire \rs2_out[20] ;
wire \rs2_out[21] ;
wire \rs2_out[22] ;
wire \rs2_out[23] ;
wire \rs2_out[24] ;
wire \rs2_out[25] ;
wire \rs2_out[26] ;
wire \rs2_out[27] ;
wire \rs2_out[28] ;
wire \rs2_out[29] ;
wire \rs2_out[30] ;
wire \rs2_out[31] ;
wire \PC_count_o[0] ;
wire \PC_count_o[1] ;
wire \PC_count_o[2] ;
wire \PC_count_o[3] ;
wire \PC_count_o[4] ;
wire \PC_count_o[5] ;
wire \PC_count_o[6] ;
wire \PC_count_o[7] ;
wire \PC_count_o[8] ;
wire \PC_count_o[9] ;
wire \PC_count_o[10] ;
wire \PC_count_o[11] ;
wire \PC_count_o[12] ;
wire \PC_count_o[13] ;
wire \PC_count_o[14] ;
wire \PC_count_o[15] ;
wire \PC_count_o[16] ;
wire \PC_count_o[17] ;
wire \PC_count_o[18] ;
wire \PC_count_o[19] ;
wire \PC_count_o[20] ;
wire \PC_count_o[21] ;
wire \PC_count_o[22] ;
wire \PC_count_o[23] ;
wire \PC_count_o[24] ;
wire \PC_count_o[25] ;
wire \PC_count_o[26] ;
wire \PC_count_o[27] ;
wire \PC_count_o[28] ;
wire \PC_count_o[29] ;
wire \PC_count_o[30] ;
wire \PC_count_o[31] ;

assign ALU_carry = ALU_overflow ;
assign ALU_carry = \imm[0] ;
assign ALU_carry = \imm[1] ;
assign ALU_carry = \imm[2] ;
assign ALU_carry = \imm[3] ;
assign ALU_carry = \imm[4] ;
assign ALU_carry = \imm[5] ;
assign ALU_carry = \imm[6] ;
assign ALU_carry = \imm[7] ;
assign ALU_carry = \imm[8] ;
assign ALU_carry = \imm[9] ;
assign ALU_carry = \imm[10] ;
assign ALU_carry = \imm[11] ;
assign ALU_carry = \imm[12] ;
assign ALU_carry = \imm[13] ;
assign ALU_carry = \imm[14] ;
assign ALU_carry = \imm[15] ;
assign ALU_carry = \imm[16] ;
assign ALU_carry = \imm[17] ;
assign ALU_carry = \imm[18] ;
assign ALU_carry = \imm[19] ;
assign ALU_carry = \imm[20] ;
assign ALU_carry = \imm[21] ;
assign ALU_carry = \imm[22] ;
assign ALU_carry = \imm[23] ;
assign ALU_carry = \imm[24] ;
assign ALU_carry = \imm[25] ;
assign ALU_carry = \imm[26] ;
assign ALU_carry = \imm[27] ;
assign ALU_carry = \imm[28] ;
assign ALU_carry = \imm[29] ;
assign ALU_carry = \imm[30] ;
assign ALU_carry = \imm[31] ;
assign ALU_carry = \rd[0] ;
assign ALU_carry = \rd[1] ;
assign ALU_carry = \rd[2] ;
assign ALU_carry = \rd[3] ;
assign ALU_carry = \rd[4] ;
assign ALU_carry = \ALU_ctrl[0] ;
assign ALU_carry = \ALU_ctrl[1] ;
assign ALU_carry = \ALU_ctrl[2] ;
assign ALU_carry = \ALU_ctrl[3] ;
assign ALU_carry = \rs1_out[0] ;
assign ALU_carry = \rs1_out[1] ;
assign ALU_carry = \rs1_out[2] ;
assign ALU_carry = \rs1_out[3] ;
assign ALU_carry = \rs1_out[4] ;
assign ALU_carry = \rs1_out[5] ;
assign ALU_carry = \rs1_out[6] ;
assign ALU_carry = \rs1_out[7] ;
assign ALU_carry = \rs1_out[8] ;
assign ALU_carry = \rs1_out[9] ;
assign ALU_carry = \rs1_out[10] ;
assign ALU_carry = \rs1_out[11] ;
assign ALU_carry = \rs1_out[12] ;
assign ALU_carry = \rs1_out[13] ;
assign ALU_carry = \rs1_out[14] ;
assign ALU_carry = \rs1_out[15] ;
assign ALU_carry = \rs1_out[16] ;
assign ALU_carry = \rs1_out[17] ;
assign ALU_carry = \rs1_out[18] ;
assign ALU_carry = \rs1_out[19] ;
assign ALU_carry = \rs1_out[20] ;
assign ALU_carry = \rs1_out[21] ;
assign ALU_carry = \rs1_out[22] ;
assign ALU_carry = \rs1_out[23] ;
assign ALU_carry = \rs1_out[24] ;
assign ALU_carry = \rs1_out[25] ;
assign ALU_carry = \rs1_out[26] ;
assign ALU_carry = \rs1_out[27] ;
assign ALU_carry = \rs1_out[28] ;
assign ALU_carry = \rs1_out[29] ;
assign ALU_carry = \rs1_out[30] ;
assign ALU_carry = \rs1_out[31] ;
assign ALU_carry = \rs2_out[0] ;
assign ALU_carry = \rs2_out[1] ;
assign ALU_carry = \rs2_out[2] ;
assign ALU_carry = \rs2_out[3] ;
assign ALU_carry = \rs2_out[4] ;
assign ALU_carry = \rs2_out[5] ;
assign ALU_carry = \rs2_out[6] ;
assign ALU_carry = \rs2_out[7] ;
assign ALU_carry = \rs2_out[8] ;
assign ALU_carry = \rs2_out[9] ;
assign ALU_carry = \rs2_out[10] ;
assign ALU_carry = \rs2_out[11] ;
assign ALU_carry = \rs2_out[12] ;
assign ALU_carry = \rs2_out[13] ;
assign ALU_carry = \rs2_out[14] ;
assign ALU_carry = \rs2_out[15] ;
assign ALU_carry = \rs2_out[16] ;
assign ALU_carry = \rs2_out[17] ;
assign ALU_carry = \rs2_out[18] ;
assign ALU_carry = \rs2_out[19] ;
assign ALU_carry = \rs2_out[20] ;
assign ALU_carry = \rs2_out[21] ;
assign ALU_carry = \rs2_out[22] ;
assign ALU_carry = \rs2_out[23] ;
assign ALU_carry = \rs2_out[24] ;
assign ALU_carry = \rs2_out[25] ;
assign ALU_carry = \rs2_out[26] ;
assign ALU_carry = \rs2_out[27] ;
assign ALU_carry = \rs2_out[28] ;
assign ALU_carry = \rs2_out[29] ;
assign ALU_carry = \rs2_out[30] ;
assign ALU_carry = \rs2_out[31] ;
assign ALU_carry = \PC_count_o[0] ;
assign ALU_carry = \PC_count_o[1] ;
assign PC_count_o[2] = \PC_count_o[2] ;
assign PC_count_o[3] = \PC_count_o[3] ;
assign PC_count_o[4] = \PC_count_o[4] ;
assign PC_count_o[5] = \PC_count_o[5] ;
assign PC_count_o[6] = \PC_count_o[6] ;
assign PC_count_o[7] = \PC_count_o[7] ;
assign PC_count_o[8] = \PC_count_o[8] ;
assign PC_count_o[9] = \PC_count_o[9] ;
assign PC_count_o[10] = \PC_count_o[10] ;
assign PC_count_o[11] = \PC_count_o[11] ;
assign PC_count_o[12] = \PC_count_o[12] ;
assign PC_count_o[13] = \PC_count_o[13] ;
assign PC_count_o[14] = \PC_count_o[14] ;
assign PC_count_o[15] = \PC_count_o[15] ;
assign PC_count_o[16] = \PC_count_o[16] ;
assign PC_count_o[17] = \PC_count_o[17] ;
assign PC_count_o[18] = \PC_count_o[18] ;
assign PC_count_o[19] = \PC_count_o[19] ;
assign PC_count_o[20] = \PC_count_o[20] ;
assign PC_count_o[21] = \PC_count_o[21] ;
assign PC_count_o[22] = \PC_count_o[22] ;
assign PC_count_o[23] = \PC_count_o[23] ;
assign PC_count_o[24] = \PC_count_o[24] ;
assign PC_count_o[25] = \PC_count_o[25] ;
assign PC_count_o[26] = \PC_count_o[26] ;
assign PC_count_o[27] = \PC_count_o[27] ;
assign PC_count_o[28] = \PC_count_o[28] ;
assign PC_count_o[29] = \PC_count_o[29] ;
assign PC_count_o[30] = \PC_count_o[30] ;
assign PC_count_o[31] = \PC_count_o[31] ;

AND2_X4 _136_ ( .A1(\PC_count_o[3] ), .A2(\PC_count_o[2] ), .ZN(_130_ ) );
AND2_X4 _137_ ( .A1(\PC_count_o[5] ), .A2(\PC_count_o[4] ), .ZN(_131_ ) );
AND2_X4 _138_ ( .A1(_130_ ), .A2(_131_ ), .ZN(_132_ ) );
AND4_X1 _139_ ( .A1(\PC_count_o[9] ), .A2(\PC_count_o[8] ), .A3(\PC_count_o[7] ), .A4(\PC_count_o[6] ), .ZN(_030_ ) );
AND2_X4 _140_ ( .A1(_132_ ), .A2(_030_ ), .ZN(_031_ ) );
INV_X1 _141_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_032_ ) );
AND2_X1 _142_ ( .A1(_031_ ), .A2(_032_ ), .ZN(_033_ ) );
INV_X1 _143_ ( .A(reset ), .ZN(_034_ ) );
OAI21_X1 _144_ ( .A(_034_ ), .B1(_031_ ), .B2(_032_ ), .ZN(_035_ ) );
NOR2_X1 _145_ ( .A1(_033_ ), .A2(_035_ ), .ZN(_000_ ) );
NAND3_X1 _146_ ( .A1(_132_ ), .A2(\PC_count_o[7] ), .A3(\PC_count_o[6] ), .ZN(_036_ ) );
NOR2_X1 _147_ ( .A1(_036_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_037_ ) );
XNOR2_X1 _148_ ( .A(_037_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_038_ ) );
CLKBUF_X2 _149_ ( .A(_034_ ), .Z(_039_ ) );
AND2_X1 _150_ ( .A1(_038_ ), .A2(_039_ ), .ZN(_001_ ) );
AND2_X4 _151_ ( .A1(\PC_count_o[13] ), .A2(\PC_count_o[12] ), .ZN(_040_ ) );
AND3_X4 _152_ ( .A1(_040_ ), .A2(\PC_count_o[11] ), .A3(\PC_count_o[10] ), .ZN(_041_ ) );
AND2_X1 _153_ ( .A1(\PC_count_o[15] ), .A2(\PC_count_o[14] ), .ZN(_042_ ) );
AND4_X4 _154_ ( .A1(\PC_count_o[16] ), .A2(_041_ ), .A3(\PC_count_o[17] ), .A4(_042_ ), .ZN(_043_ ) );
AND2_X4 _155_ ( .A1(_043_ ), .A2(_031_ ), .ZN(_044_ ) );
AND4_X1 _156_ ( .A1(\PC_count_o[24] ), .A2(\PC_count_o[23] ), .A3(\PC_count_o[25] ), .A4(\PC_count_o[22] ), .ZN(_045_ ) );
AND2_X1 _157_ ( .A1(\PC_count_o[19] ), .A2(\PC_count_o[18] ), .ZN(_046_ ) );
AND4_X1 _158_ ( .A1(\PC_count_o[20] ), .A2(_045_ ), .A3(\PC_count_o[21] ), .A4(_046_ ), .ZN(_047_ ) );
AND2_X4 _159_ ( .A1(_044_ ), .A2(_047_ ), .ZN(_048_ ) );
NAND3_X4 _160_ ( .A1(_048_ ), .A2(\PC_count_o[27] ), .A3(\PC_count_o[26] ), .ZN(_049_ ) );
OR3_X4 _161_ ( .A1(_049_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_050_ ) );
OAI21_X1 _162_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_049_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_051_ ) );
AND3_X1 _163_ ( .A1(_050_ ), .A2(_039_ ), .A3(_051_ ), .ZN(_002_ ) );
NOR2_X1 _164_ ( .A1(_049_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_052_ ) );
INV_X1 _165_ ( .A(_052_ ), .ZN(_053_ ) );
AOI21_X1 _166_ ( .A(reset ), .B1(_049_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_054_ ) );
AND2_X1 _167_ ( .A1(_053_ ), .A2(_054_ ), .ZN(_003_ ) );
INV_X1 _168_ ( .A(_048_ ), .ZN(_055_ ) );
OR3_X4 _169_ ( .A1(_055_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_056_ ) );
OAI21_X1 _170_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_055_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_057_ ) );
AND3_X1 _171_ ( .A1(_056_ ), .A2(_039_ ), .A3(_057_ ), .ZN(_004_ ) );
NOR2_X1 _172_ ( .A1(_055_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_058_ ) );
INV_X1 _173_ ( .A(_058_ ), .ZN(_059_ ) );
AOI21_X1 _174_ ( .A(reset ), .B1(_055_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_060_ ) );
AND2_X1 _175_ ( .A1(_059_ ), .A2(_060_ ), .ZN(_005_ ) );
AND3_X1 _176_ ( .A1(_046_ ), .A2(\PC_count_o[20] ), .A3(\PC_count_o[21] ), .ZN(_061_ ) );
AND3_X4 _177_ ( .A1(_043_ ), .A2(_031_ ), .A3(_061_ ), .ZN(_062_ ) );
AND3_X4 _178_ ( .A1(_062_ ), .A2(\PC_count_o[23] ), .A3(\PC_count_o[22] ), .ZN(_063_ ) );
INV_X2 _179_ ( .A(_063_ ), .ZN(_064_ ) );
OR3_X4 _180_ ( .A1(_064_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_065_ ) );
OAI21_X1 _181_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_064_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_066_ ) );
AND3_X1 _182_ ( .A1(_065_ ), .A2(_039_ ), .A3(_066_ ), .ZN(_006_ ) );
NOR2_X1 _183_ ( .A1(_064_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_067_ ) );
INV_X1 _184_ ( .A(_067_ ), .ZN(_068_ ) );
AOI21_X1 _185_ ( .A(reset ), .B1(_064_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_069_ ) );
AND2_X1 _186_ ( .A1(_068_ ), .A2(_069_ ), .ZN(_007_ ) );
INV_X1 _187_ ( .A(_062_ ), .ZN(_070_ ) );
OR3_X1 _188_ ( .A1(_070_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_071_ ) );
OAI21_X1 _189_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_070_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_072_ ) );
AND3_X1 _190_ ( .A1(_071_ ), .A2(_039_ ), .A3(_072_ ), .ZN(_008_ ) );
NOR2_X1 _191_ ( .A1(_070_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_073_ ) );
INV_X1 _192_ ( .A(_073_ ), .ZN(_074_ ) );
AOI21_X1 _193_ ( .A(reset ), .B1(_070_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_075_ ) );
AND2_X1 _194_ ( .A1(_074_ ), .A2(_075_ ), .ZN(_009_ ) );
NAND3_X1 _195_ ( .A1(_043_ ), .A2(_031_ ), .A3(_046_ ), .ZN(_076_ ) );
OR3_X1 _196_ ( .A1(_076_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_077_ ) );
OAI21_X1 _197_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_076_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_078_ ) );
AND3_X1 _198_ ( .A1(_077_ ), .A2(_039_ ), .A3(_078_ ), .ZN(_010_ ) );
NOR2_X1 _199_ ( .A1(_076_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_079_ ) );
INV_X1 _200_ ( .A(_079_ ), .ZN(_080_ ) );
AOI21_X1 _201_ ( .A(reset ), .B1(_076_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_081_ ) );
AND2_X1 _202_ ( .A1(_080_ ), .A2(_081_ ), .ZN(_011_ ) );
INV_X1 _203_ ( .A(_037_ ), .ZN(_082_ ) );
AOI21_X1 _204_ ( .A(reset ), .B1(_036_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_083_ ) );
AND2_X1 _205_ ( .A1(_082_ ), .A2(_083_ ), .ZN(_012_ ) );
INV_X1 _206_ ( .A(_044_ ), .ZN(_084_ ) );
OR3_X1 _207_ ( .A1(_084_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_085_ ) );
OAI21_X1 _208_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_084_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_086_ ) );
AND3_X1 _209_ ( .A1(_085_ ), .A2(_039_ ), .A3(_086_ ), .ZN(_013_ ) );
NOR2_X1 _210_ ( .A1(_084_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_087_ ) );
INV_X1 _211_ ( .A(_087_ ), .ZN(_088_ ) );
AOI21_X1 _212_ ( .A(reset ), .B1(_084_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_089_ ) );
AND2_X1 _213_ ( .A1(_088_ ), .A2(_089_ ), .ZN(_014_ ) );
AND3_X1 _214_ ( .A1(_031_ ), .A2(_041_ ), .A3(_042_ ), .ZN(_090_ ) );
INV_X1 _215_ ( .A(_090_ ), .ZN(_091_ ) );
OR3_X1 _216_ ( .A1(_091_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_092_ ) );
OAI21_X1 _217_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_091_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_093_ ) );
AND3_X1 _218_ ( .A1(_092_ ), .A2(_039_ ), .A3(_093_ ), .ZN(_015_ ) );
AND3_X1 _219_ ( .A1(_031_ ), .A2(\PC_count_o[11] ), .A3(\PC_count_o[10] ), .ZN(_094_ ) );
NAND3_X1 _220_ ( .A1(_094_ ), .A2(_040_ ), .A3(_042_ ), .ZN(_095_ ) );
OR2_X1 _221_ ( .A1(_095_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_096_ ) );
AOI21_X1 _222_ ( .A(reset ), .B1(_091_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_097_ ) );
AND2_X1 _223_ ( .A1(_096_ ), .A2(_097_ ), .ZN(_016_ ) );
AND3_X1 _224_ ( .A1(_041_ ), .A2(_132_ ), .A3(_030_ ), .ZN(_098_ ) );
INV_X1 _225_ ( .A(_098_ ), .ZN(_099_ ) );
OR3_X1 _226_ ( .A1(_099_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_100_ ) );
OAI21_X1 _227_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_099_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_101_ ) );
AND3_X1 _228_ ( .A1(_100_ ), .A2(_034_ ), .A3(_101_ ), .ZN(_017_ ) );
NAND2_X1 _229_ ( .A1(_094_ ), .A2(_040_ ), .ZN(_102_ ) );
OR2_X1 _230_ ( .A1(_102_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_103_ ) );
AOI21_X1 _231_ ( .A(reset ), .B1(_099_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_104_ ) );
AND2_X1 _232_ ( .A1(_103_ ), .A2(_104_ ), .ZN(_018_ ) );
INV_X1 _233_ ( .A(_094_ ), .ZN(_105_ ) );
OR3_X1 _234_ ( .A1(_105_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_106_ ) );
OAI21_X1 _235_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ), .B1(_105_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_107_ ) );
AND3_X1 _236_ ( .A1(_106_ ), .A2(_034_ ), .A3(_107_ ), .ZN(_019_ ) );
NOR2_X1 _237_ ( .A1(_105_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_108_ ) );
INV_X1 _238_ ( .A(_108_ ), .ZN(_109_ ) );
AOI21_X1 _239_ ( .A(reset ), .B1(_105_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_110_ ) );
AND2_X1 _240_ ( .A1(_109_ ), .A2(_110_ ), .ZN(_020_ ) );
INV_X1 _241_ ( .A(_033_ ), .ZN(_111_ ) );
AOI21_X1 _242_ ( .A(reset ), .B1(_111_ ), .B2(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_112_ ) );
INV_X1 _243_ ( .A(_031_ ), .ZN(_113_ ) );
OR3_X1 _244_ ( .A1(_113_ ), .A2(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_B_$_XOR__Y_B ), .A3(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_114_ ) );
AND2_X1 _245_ ( .A1(_112_ ), .A2(_114_ ), .ZN(_021_ ) );
INV_X1 _246_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_115_ ) );
AND2_X1 _247_ ( .A1(_132_ ), .A2(_115_ ), .ZN(_116_ ) );
XNOR2_X1 _248_ ( .A(_116_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_117_ ) );
AND2_X1 _249_ ( .A1(_117_ ), .A2(_039_ ), .ZN(_022_ ) );
OAI21_X1 _250_ ( .A(_034_ ), .B1(_132_ ), .B2(_115_ ), .ZN(_118_ ) );
NOR2_X1 _251_ ( .A1(_116_ ), .A2(_118_ ), .ZN(_023_ ) );
INV_X1 _252_ ( .A(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_119_ ) );
AND2_X1 _253_ ( .A1(_130_ ), .A2(_119_ ), .ZN(_120_ ) );
XNOR2_X1 _254_ ( .A(_120_ ), .B(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ), .ZN(_121_ ) );
AND2_X1 _255_ ( .A1(_121_ ), .A2(_039_ ), .ZN(_024_ ) );
OAI21_X1 _256_ ( .A(_034_ ), .B1(_130_ ), .B2(_119_ ), .ZN(_122_ ) );
NOR2_X1 _257_ ( .A1(_120_ ), .A2(_122_ ), .ZN(_025_ ) );
NOR2_X1 _258_ ( .A1(\PC_count_o[3] ), .A2(\PC_count_o[2] ), .ZN(_123_ ) );
NOR3_X1 _259_ ( .A1(_130_ ), .A2(_123_ ), .A3(reset ), .ZN(_026_ ) );
NOR2_X1 _260_ ( .A1(reset ), .A2(\PC_count_o[2] ), .ZN(_027_ ) );
AND4_X1 _261_ ( .A1(\PC_count_o[29] ), .A2(\PC_count_o[28] ), .A3(\PC_count_o[27] ), .A4(\PC_count_o[26] ), .ZN(_124_ ) );
NAND3_X1 _262_ ( .A1(_044_ ), .A2(_047_ ), .A3(_124_ ), .ZN(_125_ ) );
NOR2_X1 _263_ ( .A1(_125_ ), .A2(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_126_ ) );
INV_X1 _264_ ( .A(_126_ ), .ZN(_127_ ) );
AOI21_X1 _265_ ( .A(reset ), .B1(_125_ ), .B2(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ), .ZN(_128_ ) );
AND2_X1 _266_ ( .A1(_127_ ), .A2(_128_ ), .ZN(_028_ ) );
AOI21_X1 _267_ ( .A(reset ), .B1(_126_ ), .B2(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_129_ ) );
OAI21_X1 _268_ ( .A(_129_ ), .B1(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_126_ ), .ZN(_029_ ) );
CLKGATE_X1 _269_ ( .CK(clk ), .E(\i0.state_$_SDFFE_PP0P__Q_E ), .GCK(_133_ ) );
CLKGATE_X1 _270_ ( .CK(clk ), .E(\i0.state_$_SDFFE_PP0P__Q_E ), .GCK(_134_ ) );
LOGIC1_X1 _271_ ( .Z(\i0.state_$_SDFFE_PP0P__Q_E ) );
LOGIC0_X1 _272_ ( .Z(ALU_carry ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q ( .D(_000_ ), .CK(_134_ ), .Q(\PC_count_o[10] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_21_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_1 ( .D(_001_ ), .CK(_134_ ), .Q(\PC_count_o[9] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_22_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_10 ( .D(_002_ ), .CK(_133_ ), .Q(\PC_count_o[29] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_2_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_11 ( .D(_003_ ), .CK(_133_ ), .Q(\PC_count_o[28] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_3_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_12 ( .D(_004_ ), .CK(_133_ ), .Q(\PC_count_o[27] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_4_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_13 ( .D(_005_ ), .CK(_133_ ), .Q(\PC_count_o[26] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_5_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_14 ( .D(_006_ ), .CK(_133_ ), .Q(\PC_count_o[25] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_6_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_15 ( .D(_007_ ), .CK(_133_ ), .Q(\PC_count_o[24] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_7_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_16 ( .D(_008_ ), .CK(_133_ ), .Q(\PC_count_o[23] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_8_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_17 ( .D(_009_ ), .CK(_133_ ), .Q(\PC_count_o[22] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_9_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_18 ( .D(_010_ ), .CK(_133_ ), .Q(\PC_count_o[21] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_10_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_19 ( .D(_011_ ), .CK(_133_ ), .Q(\PC_count_o[20] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_11_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_2 ( .D(_012_ ), .CK(_134_ ), .Q(\PC_count_o[8] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_23_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_20 ( .D(_013_ ), .CK(_133_ ), .Q(\PC_count_o[19] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_12_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_21 ( .D(_014_ ), .CK(_133_ ), .Q(\PC_count_o[18] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_13_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_22 ( .D(_015_ ), .CK(_133_ ), .Q(\PC_count_o[17] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_14_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_23 ( .D(_016_ ), .CK(_133_ ), .Q(\PC_count_o[16] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_15_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_24 ( .D(_017_ ), .CK(_133_ ), .Q(\PC_count_o[15] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_16_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_25 ( .D(_018_ ), .CK(_133_ ), .Q(\PC_count_o[14] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_17_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_26 ( .D(_019_ ), .CK(_133_ ), .Q(\PC_count_o[13] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_18_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_27 ( .D(_020_ ), .CK(_133_ ), .Q(\PC_count_o[12] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_28 ( .D(_021_ ), .CK(_133_ ), .Q(\PC_count_o[11] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_20_B_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_3 ( .D(_022_ ), .CK(_134_ ), .Q(\PC_count_o[7] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_24_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_4 ( .D(_023_ ), .CK(_134_ ), .Q(\PC_count_o[6] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_25_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_5 ( .D(_024_ ), .CK(_134_ ), .Q(\PC_count_o[5] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_26_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_6 ( .D(_025_ ), .CK(_134_ ), .Q(\PC_count_o[4] ), .QN(\i7._io_pc_next_T_26_$_ANDNOT__Y_27_B_$_OR__Y_A_$_MUX__Y_B_$_XOR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_7 ( .D(_026_ ), .CK(_134_ ), .Q(\PC_count_o[3] ), .QN(_135_ ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_8 ( .D(_027_ ), .CK(_134_ ), .Q(\PC_count_o[2] ), .QN(ALU_carry_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ANDNOT__Y_A_$_NAND__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \i0.state_$_SDFFE_PP0P__Q_9 ( .D(_028_ ), .CK(_133_ ), .Q(\PC_count_o[30] ), .QN(ALU_overflow_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B ) );
DFF_X1 \i0.state_$_SDFFE_PP1P__Q ( .D(_029_ ), .CK(_133_ ), .Q(\PC_count_o[31] ), .QN(ALU_overflow_$_ANDNOT__Y_A_$_OR__Y_B ) );

endmodule
